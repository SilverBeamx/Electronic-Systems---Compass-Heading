library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.numeric_std.all;

entity atan_lut_4096_8bit is
  port (
    address  : in  std_logic_vector(11 downto 0);
    atan_out : out std_logic_vector(7 downto 0)
  );
end entity;

architecture rtl of atan_lut_4096_8bit is

  type LUT_t is array (natural range 0 to 4095) of natural;
  constant LUT: LUT_t := (
    0 => 0,               -- (000000.000000 | 0.0)          => (000.00000 | 0.0)             
    1 => 0,               -- (000000.000001 | 0.015625)     => (000.00000 | 0.0)             
    2 => 0,               -- (000000.000010 | 0.03125)      => (000.00000 | 0.0)             
    3 => 1,               -- (000000.000011 | 0.046875)     => (000.00001 | 0.03125)         
    4 => 1,               -- (000000.000100 | 0.0625)       => (000.00001 | 0.03125)         
    5 => 2,               -- (000000.000101 | 0.078125)     => (000.00010 | 0.0625)          
    6 => 2,               -- (000000.000110 | 0.09375)      => (000.00010 | 0.0625)          
    7 => 3,               -- (000000.000111 | 0.109375)     => (000.00011 | 0.09375)         
    8 => 3,               -- (000000.001000 | 0.125)        => (000.00011 | 0.09375)         
    9 => 4,               -- (000000.001001 | 0.140625)     => (000.00100 | 0.125)           
    10 => 4,              -- (000000.001010 | 0.15625)      => (000.00100 | 0.125)           
    11 => 5,              -- (000000.001011 | 0.171875)     => (000.00101 | 0.15625)         
    12 => 5,              -- (000000.001100 | 0.1875)       => (000.00101 | 0.15625)         
    13 => 6,              -- (000000.001101 | 0.203125)     => (000.00110 | 0.1875)          
    14 => 6,              -- (000000.001110 | 0.21875)      => (000.00110 | 0.1875)          
    15 => 7,              -- (000000.001111 | 0.234375)     => (000.00111 | 0.21875)         
    16 => 7,              -- (000000.010000 | 0.25)         => (000.00111 | 0.21875)         
    17 => 8,              -- (000000.010001 | 0.265625)     => (000.01000 | 0.25)            
    18 => 8,              -- (000000.010010 | 0.28125)      => (000.01000 | 0.25)            
    19 => 9,              -- (000000.010011 | 0.296875)     => (000.01001 | 0.28125)         
    20 => 9,              -- (000000.010100 | 0.3125)       => (000.01001 | 0.28125)         
    21 => 10,             -- (000000.010101 | 0.328125)     => (000.01010 | 0.3125)          
    22 => 10,             -- (000000.010110 | 0.34375)      => (000.01010 | 0.3125)          
    23 => 11,             -- (000000.010111 | 0.359375)     => (000.01011 | 0.34375)         
    24 => 11,             -- (000000.011000 | 0.375)        => (000.01011 | 0.34375)         
    25 => 11,             -- (000000.011001 | 0.390625)     => (000.01011 | 0.34375)         
    26 => 12,             -- (000000.011010 | 0.40625)      => (000.01100 | 0.375)           
    27 => 12,             -- (000000.011011 | 0.421875)     => (000.01100 | 0.375)           
    28 => 13,             -- (000000.011100 | 0.4375)       => (000.01101 | 0.40625)         
    29 => 13,             -- (000000.011101 | 0.453125)     => (000.01101 | 0.40625)         
    30 => 14,             -- (000000.011110 | 0.46875)      => (000.01110 | 0.4375)          
    31 => 14,             -- (000000.011111 | 0.484375)     => (000.01110 | 0.4375)          
    32 => 14,             -- (000000.100000 | 0.5)          => (000.01110 | 0.4375)          
    33 => 15,             -- (000000.100001 | 0.515625)     => (000.01111 | 0.46875)         
    34 => 15,             -- (000000.100010 | 0.53125)      => (000.01111 | 0.46875)         
    35 => 16,             -- (000000.100011 | 0.546875)     => (000.10000 | 0.5)             
    36 => 16,             -- (000000.100100 | 0.5625)       => (000.10000 | 0.5)             
    37 => 16,             -- (000000.100101 | 0.578125)     => (000.10000 | 0.5)             
    38 => 17,             -- (000000.100110 | 0.59375)      => (000.10001 | 0.53125)         
    39 => 17,             -- (000000.100111 | 0.609375)     => (000.10001 | 0.53125)         
    40 => 17,             -- (000000.101000 | 0.625)        => (000.10001 | 0.53125)         
    41 => 18,             -- (000000.101001 | 0.640625)     => (000.10010 | 0.5625)          
    42 => 18,             -- (000000.101010 | 0.65625)      => (000.10010 | 0.5625)          
    43 => 18,             -- (000000.101011 | 0.671875)     => (000.10010 | 0.5625)          
    44 => 19,             -- (000000.101100 | 0.6875)       => (000.10011 | 0.59375)         
    45 => 19,             -- (000000.101101 | 0.703125)     => (000.10011 | 0.59375)         
    46 => 19,             -- (000000.101110 | 0.71875)      => (000.10011 | 0.59375)         
    47 => 20,             -- (000000.101111 | 0.734375)     => (000.10100 | 0.625)           
    48 => 20,             -- (000000.110000 | 0.75)         => (000.10100 | 0.625)           
    49 => 20,             -- (000000.110001 | 0.765625)     => (000.10100 | 0.625)           
    50 => 21,             -- (000000.110010 | 0.78125)      => (000.10101 | 0.65625)         
    51 => 21,             -- (000000.110011 | 0.796875)     => (000.10101 | 0.65625)         
    52 => 21,             -- (000000.110100 | 0.8125)       => (000.10101 | 0.65625)         
    53 => 22,             -- (000000.110101 | 0.828125)     => (000.10110 | 0.6875)          
    54 => 22,             -- (000000.110110 | 0.84375)      => (000.10110 | 0.6875)          
    55 => 22,             -- (000000.110111 | 0.859375)     => (000.10110 | 0.6875)          
    56 => 23,             -- (000000.111000 | 0.875)        => (000.10111 | 0.71875)         
    57 => 23,             -- (000000.111001 | 0.890625)     => (000.10111 | 0.71875)         
    58 => 23,             -- (000000.111010 | 0.90625)      => (000.10111 | 0.71875)         
    59 => 23,             -- (000000.111011 | 0.921875)     => (000.10111 | 0.71875)         
    60 => 24,             -- (000000.111100 | 0.9375)       => (000.11000 | 0.75)            
    61 => 24,             -- (000000.111101 | 0.953125)     => (000.11000 | 0.75)            
    62 => 24,             -- (000000.111110 | 0.96875)      => (000.11000 | 0.75)            
    63 => 24,             -- (000000.111111 | 0.984375)     => (000.11000 | 0.75)            
    64 => 25,             -- (000001.000000 | 1.0)          => (000.11001 | 0.78125)         
    65 => 25,             -- (000001.000001 | 1.015625)     => (000.11001 | 0.78125)         
    66 => 25,             -- (000001.000010 | 1.03125)      => (000.11001 | 0.78125)         
    67 => 25,             -- (000001.000011 | 1.046875)     => (000.11001 | 0.78125)         
    68 => 26,             -- (000001.000100 | 1.0625)       => (000.11010 | 0.8125)          
    69 => 26,             -- (000001.000101 | 1.078125)     => (000.11010 | 0.8125)          
    70 => 26,             -- (000001.000110 | 1.09375)      => (000.11010 | 0.8125)          
    71 => 26,             -- (000001.000111 | 1.109375)     => (000.11010 | 0.8125)          
    72 => 27,             -- (000001.001000 | 1.125)        => (000.11011 | 0.84375)         
    73 => 27,             -- (000001.001001 | 1.140625)     => (000.11011 | 0.84375)         
    74 => 27,             -- (000001.001010 | 1.15625)      => (000.11011 | 0.84375)         
    75 => 27,             -- (000001.001011 | 1.171875)     => (000.11011 | 0.84375)         
    76 => 27,             -- (000001.001100 | 1.1875)       => (000.11011 | 0.84375)         
    77 => 28,             -- (000001.001101 | 1.203125)     => (000.11100 | 0.875)           
    78 => 28,             -- (000001.001110 | 1.21875)      => (000.11100 | 0.875)           
    79 => 28,             -- (000001.001111 | 1.234375)     => (000.11100 | 0.875)           
    80 => 28,             -- (000001.010000 | 1.25)         => (000.11100 | 0.875)           
    81 => 28,             -- (000001.010001 | 1.265625)     => (000.11100 | 0.875)           
    82 => 29,             -- (000001.010010 | 1.28125)      => (000.11101 | 0.90625)         
    83 => 29,             -- (000001.010011 | 1.296875)     => (000.11101 | 0.90625)         
    84 => 29,             -- (000001.010100 | 1.3125)       => (000.11101 | 0.90625)         
    85 => 29,             -- (000001.010101 | 1.328125)     => (000.11101 | 0.90625)         
    86 => 29,             -- (000001.010110 | 1.34375)      => (000.11101 | 0.90625)         
    87 => 29,             -- (000001.010111 | 1.359375)     => (000.11101 | 0.90625)         
    88 => 30,             -- (000001.011000 | 1.375)        => (000.11110 | 0.9375)          
    89 => 30,             -- (000001.011001 | 1.390625)     => (000.11110 | 0.9375)          
    90 => 30,             -- (000001.011010 | 1.40625)      => (000.11110 | 0.9375)          
    91 => 30,             -- (000001.011011 | 1.421875)     => (000.11110 | 0.9375)          
    92 => 30,             -- (000001.011100 | 1.4375)       => (000.11110 | 0.9375)          
    93 => 30,             -- (000001.011101 | 1.453125)     => (000.11110 | 0.9375)          
    94 => 31,             -- (000001.011110 | 1.46875)      => (000.11111 | 0.96875)         
    95 => 31,             -- (000001.011111 | 1.484375)     => (000.11111 | 0.96875)         
    96 => 31,             -- (000001.100000 | 1.5)          => (000.11111 | 0.96875)         
    97 => 31,             -- (000001.100001 | 1.515625)     => (000.11111 | 0.96875)         
    98 => 31,             -- (000001.100010 | 1.53125)      => (000.11111 | 0.96875)         
    99 => 31,             -- (000001.100011 | 1.546875)     => (000.11111 | 0.96875)         
    100 => 32,            -- (000001.100100 | 1.5625)       => (001.00000 | 1.0)             
    101 => 32,            -- (000001.100101 | 1.578125)     => (001.00000 | 1.0)             
    102 => 32,            -- (000001.100110 | 1.59375)      => (001.00000 | 1.0)             
    103 => 32,            -- (000001.100111 | 1.609375)     => (001.00000 | 1.0)             
    104 => 32,            -- (000001.101000 | 1.625)        => (001.00000 | 1.0)             
    105 => 32,            -- (000001.101001 | 1.640625)     => (001.00000 | 1.0)             
    106 => 32,            -- (000001.101010 | 1.65625)      => (001.00000 | 1.0)             
    107 => 33,            -- (000001.101011 | 1.671875)     => (001.00001 | 1.03125)         
    108 => 33,            -- (000001.101100 | 1.6875)       => (001.00001 | 1.03125)         
    109 => 33,            -- (000001.101101 | 1.703125)     => (001.00001 | 1.03125)         
    110 => 33,            -- (000001.101110 | 1.71875)      => (001.00001 | 1.03125)         
    111 => 33,            -- (000001.101111 | 1.734375)     => (001.00001 | 1.03125)         
    112 => 33,            -- (000001.110000 | 1.75)         => (001.00001 | 1.03125)         
    113 => 33,            -- (000001.110001 | 1.765625)     => (001.00001 | 1.03125)         
    114 => 33,            -- (000001.110010 | 1.78125)      => (001.00001 | 1.03125)         
    115 => 34,            -- (000001.110011 | 1.796875)     => (001.00010 | 1.0625)          
    116 => 34,            -- (000001.110100 | 1.8125)       => (001.00010 | 1.0625)          
    117 => 34,            -- (000001.110101 | 1.828125)     => (001.00010 | 1.0625)          
    118 => 34,            -- (000001.110110 | 1.84375)      => (001.00010 | 1.0625)          
    119 => 34,            -- (000001.110111 | 1.859375)     => (001.00010 | 1.0625)          
    120 => 34,            -- (000001.111000 | 1.875)        => (001.00010 | 1.0625)          
    121 => 34,            -- (000001.111001 | 1.890625)     => (001.00010 | 1.0625)          
    122 => 34,            -- (000001.111010 | 1.90625)      => (001.00010 | 1.0625)          
    123 => 34,            -- (000001.111011 | 1.921875)     => (001.00010 | 1.0625)          
    124 => 35,            -- (000001.111100 | 1.9375)       => (001.00011 | 1.09375)         
    125 => 35,            -- (000001.111101 | 1.953125)     => (001.00011 | 1.09375)         
    126 => 35,            -- (000001.111110 | 1.96875)      => (001.00011 | 1.09375)         
    127 => 35,            -- (000001.111111 | 1.984375)     => (001.00011 | 1.09375)         
    128 => 35,            -- (000010.000000 | 2.0)          => (001.00011 | 1.09375)         
    129 => 35,            -- (000010.000001 | 2.015625)     => (001.00011 | 1.09375)         
    130 => 35,            -- (000010.000010 | 2.03125)      => (001.00011 | 1.09375)         
    131 => 35,            -- (000010.000011 | 2.046875)     => (001.00011 | 1.09375)         
    132 => 35,            -- (000010.000100 | 2.0625)       => (001.00011 | 1.09375)         
    133 => 35,            -- (000010.000101 | 2.078125)     => (001.00011 | 1.09375)         
    134 => 36,            -- (000010.000110 | 2.09375)      => (001.00100 | 1.125)           
    135 => 36,            -- (000010.000111 | 2.109375)     => (001.00100 | 1.125)           
    136 => 36,            -- (000010.001000 | 2.125)        => (001.00100 | 1.125)           
    137 => 36,            -- (000010.001001 | 2.140625)     => (001.00100 | 1.125)           
    138 => 36,            -- (000010.001010 | 2.15625)      => (001.00100 | 1.125)           
    139 => 36,            -- (000010.001011 | 2.171875)     => (001.00100 | 1.125)           
    140 => 36,            -- (000010.001100 | 2.1875)       => (001.00100 | 1.125)           
    141 => 36,            -- (000010.001101 | 2.203125)     => (001.00100 | 1.125)           
    142 => 36,            -- (000010.001110 | 2.21875)      => (001.00100 | 1.125)           
    143 => 36,            -- (000010.001111 | 2.234375)     => (001.00100 | 1.125)           
    144 => 36,            -- (000010.010000 | 2.25)         => (001.00100 | 1.125)           
    145 => 36,            -- (000010.010001 | 2.265625)     => (001.00100 | 1.125)           
    146 => 37,            -- (000010.010010 | 2.28125)      => (001.00101 | 1.15625)         
    147 => 37,            -- (000010.010011 | 2.296875)     => (001.00101 | 1.15625)         
    148 => 37,            -- (000010.010100 | 2.3125)       => (001.00101 | 1.15625)         
    149 => 37,            -- (000010.010101 | 2.328125)     => (001.00101 | 1.15625)         
    150 => 37,            -- (000010.010110 | 2.34375)      => (001.00101 | 1.15625)         
    151 => 37,            -- (000010.010111 | 2.359375)     => (001.00101 | 1.15625)         
    152 => 37,            -- (000010.011000 | 2.375)        => (001.00101 | 1.15625)         
    153 => 37,            -- (000010.011001 | 2.390625)     => (001.00101 | 1.15625)         
    154 => 37,            -- (000010.011010 | 2.40625)      => (001.00101 | 1.15625)         
    155 => 37,            -- (000010.011011 | 2.421875)     => (001.00101 | 1.15625)         
    156 => 37,            -- (000010.011100 | 2.4375)       => (001.00101 | 1.15625)         
    157 => 37,            -- (000010.011101 | 2.453125)     => (001.00101 | 1.15625)         
    158 => 37,            -- (000010.011110 | 2.46875)      => (001.00101 | 1.15625)         
    159 => 38,            -- (000010.011111 | 2.484375)     => (001.00110 | 1.1875)          
    160 => 38,            -- (000010.100000 | 2.5)          => (001.00110 | 1.1875)          
    161 => 38,            -- (000010.100001 | 2.515625)     => (001.00110 | 1.1875)          
    162 => 38,            -- (000010.100010 | 2.53125)      => (001.00110 | 1.1875)          
    163 => 38,            -- (000010.100011 | 2.546875)     => (001.00110 | 1.1875)          
    164 => 38,            -- (000010.100100 | 2.5625)       => (001.00110 | 1.1875)          
    165 => 38,            -- (000010.100101 | 2.578125)     => (001.00110 | 1.1875)          
    166 => 38,            -- (000010.100110 | 2.59375)      => (001.00110 | 1.1875)          
    167 => 38,            -- (000010.100111 | 2.609375)     => (001.00110 | 1.1875)          
    168 => 38,            -- (000010.101000 | 2.625)        => (001.00110 | 1.1875)          
    169 => 38,            -- (000010.101001 | 2.640625)     => (001.00110 | 1.1875)          
    170 => 38,            -- (000010.101010 | 2.65625)      => (001.00110 | 1.1875)          
    171 => 38,            -- (000010.101011 | 2.671875)     => (001.00110 | 1.1875)          
    172 => 38,            -- (000010.101100 | 2.6875)       => (001.00110 | 1.1875)          
    173 => 38,            -- (000010.101101 | 2.703125)     => (001.00110 | 1.1875)          
    174 => 38,            -- (000010.101110 | 2.71875)      => (001.00110 | 1.1875)          
    175 => 39,            -- (000010.101111 | 2.734375)     => (001.00111 | 1.21875)         
    176 => 39,            -- (000010.110000 | 2.75)         => (001.00111 | 1.21875)         
    177 => 39,            -- (000010.110001 | 2.765625)     => (001.00111 | 1.21875)         
    178 => 39,            -- (000010.110010 | 2.78125)      => (001.00111 | 1.21875)         
    179 => 39,            -- (000010.110011 | 2.796875)     => (001.00111 | 1.21875)         
    180 => 39,            -- (000010.110100 | 2.8125)       => (001.00111 | 1.21875)         
    181 => 39,            -- (000010.110101 | 2.828125)     => (001.00111 | 1.21875)         
    182 => 39,            -- (000010.110110 | 2.84375)      => (001.00111 | 1.21875)         
    183 => 39,            -- (000010.110111 | 2.859375)     => (001.00111 | 1.21875)         
    184 => 39,            -- (000010.111000 | 2.875)        => (001.00111 | 1.21875)         
    185 => 39,            -- (000010.111001 | 2.890625)     => (001.00111 | 1.21875)         
    186 => 39,            -- (000010.111010 | 2.90625)      => (001.00111 | 1.21875)         
    187 => 39,            -- (000010.111011 | 2.921875)     => (001.00111 | 1.21875)         
    188 => 39,            -- (000010.111100 | 2.9375)       => (001.00111 | 1.21875)         
    189 => 39,            -- (000010.111101 | 2.953125)     => (001.00111 | 1.21875)         
    190 => 39,            -- (000010.111110 | 2.96875)      => (001.00111 | 1.21875)         
    191 => 39,            -- (000010.111111 | 2.984375)     => (001.00111 | 1.21875)         
    192 => 39,            -- (000011.000000 | 3.0)          => (001.00111 | 1.21875)         
    193 => 40,            -- (000011.000001 | 3.015625)     => (001.01000 | 1.25)            
    194 => 40,            -- (000011.000010 | 3.03125)      => (001.01000 | 1.25)            
    195 => 40,            -- (000011.000011 | 3.046875)     => (001.01000 | 1.25)            
    196 => 40,            -- (000011.000100 | 3.0625)       => (001.01000 | 1.25)            
    197 => 40,            -- (000011.000101 | 3.078125)     => (001.01000 | 1.25)            
    198 => 40,            -- (000011.000110 | 3.09375)      => (001.01000 | 1.25)            
    199 => 40,            -- (000011.000111 | 3.109375)     => (001.01000 | 1.25)            
    200 => 40,            -- (000011.001000 | 3.125)        => (001.01000 | 1.25)            
    201 => 40,            -- (000011.001001 | 3.140625)     => (001.01000 | 1.25)            
    202 => 40,            -- (000011.001010 | 3.15625)      => (001.01000 | 1.25)            
    203 => 40,            -- (000011.001011 | 3.171875)     => (001.01000 | 1.25)            
    204 => 40,            -- (000011.001100 | 3.1875)       => (001.01000 | 1.25)            
    205 => 40,            -- (000011.001101 | 3.203125)     => (001.01000 | 1.25)            
    206 => 40,            -- (000011.001110 | 3.21875)      => (001.01000 | 1.25)            
    207 => 40,            -- (000011.001111 | 3.234375)     => (001.01000 | 1.25)            
    208 => 40,            -- (000011.010000 | 3.25)         => (001.01000 | 1.25)            
    209 => 40,            -- (000011.010001 | 3.265625)     => (001.01000 | 1.25)            
    210 => 40,            -- (000011.010010 | 3.28125)      => (001.01000 | 1.25)            
    211 => 40,            -- (000011.010011 | 3.296875)     => (001.01000 | 1.25)            
    212 => 40,            -- (000011.010100 | 3.3125)       => (001.01000 | 1.25)            
    213 => 40,            -- (000011.010101 | 3.328125)     => (001.01000 | 1.25)            
    214 => 40,            -- (000011.010110 | 3.34375)      => (001.01000 | 1.25)            
    215 => 41,            -- (000011.010111 | 3.359375)     => (001.01001 | 1.28125)         
    216 => 41,            -- (000011.011000 | 3.375)        => (001.01001 | 1.28125)         
    217 => 41,            -- (000011.011001 | 3.390625)     => (001.01001 | 1.28125)         
    218 => 41,            -- (000011.011010 | 3.40625)      => (001.01001 | 1.28125)         
    219 => 41,            -- (000011.011011 | 3.421875)     => (001.01001 | 1.28125)         
    220 => 41,            -- (000011.011100 | 3.4375)       => (001.01001 | 1.28125)         
    221 => 41,            -- (000011.011101 | 3.453125)     => (001.01001 | 1.28125)         
    222 => 41,            -- (000011.011110 | 3.46875)      => (001.01001 | 1.28125)         
    223 => 41,            -- (000011.011111 | 3.484375)     => (001.01001 | 1.28125)         
    224 => 41,            -- (000011.100000 | 3.5)          => (001.01001 | 1.28125)         
    225 => 41,            -- (000011.100001 | 3.515625)     => (001.01001 | 1.28125)         
    226 => 41,            -- (000011.100010 | 3.53125)      => (001.01001 | 1.28125)         
    227 => 41,            -- (000011.100011 | 3.546875)     => (001.01001 | 1.28125)         
    228 => 41,            -- (000011.100100 | 3.5625)       => (001.01001 | 1.28125)         
    229 => 41,            -- (000011.100101 | 3.578125)     => (001.01001 | 1.28125)         
    230 => 41,            -- (000011.100110 | 3.59375)      => (001.01001 | 1.28125)         
    231 => 41,            -- (000011.100111 | 3.609375)     => (001.01001 | 1.28125)         
    232 => 41,            -- (000011.101000 | 3.625)        => (001.01001 | 1.28125)         
    233 => 41,            -- (000011.101001 | 3.640625)     => (001.01001 | 1.28125)         
    234 => 41,            -- (000011.101010 | 3.65625)      => (001.01001 | 1.28125)         
    235 => 41,            -- (000011.101011 | 3.671875)     => (001.01001 | 1.28125)         
    236 => 41,            -- (000011.101100 | 3.6875)       => (001.01001 | 1.28125)         
    237 => 41,            -- (000011.101101 | 3.703125)     => (001.01001 | 1.28125)         
    238 => 41,            -- (000011.101110 | 3.71875)      => (001.01001 | 1.28125)         
    239 => 41,            -- (000011.101111 | 3.734375)     => (001.01001 | 1.28125)         
    240 => 41,            -- (000011.110000 | 3.75)         => (001.01001 | 1.28125)         
    241 => 41,            -- (000011.110001 | 3.765625)     => (001.01001 | 1.28125)         
    242 => 41,            -- (000011.110010 | 3.78125)      => (001.01001 | 1.28125)         
    243 => 42,            -- (000011.110011 | 3.796875)     => (001.01010 | 1.3125)          
    244 => 42,            -- (000011.110100 | 3.8125)       => (001.01010 | 1.3125)          
    245 => 42,            -- (000011.110101 | 3.828125)     => (001.01010 | 1.3125)          
    246 => 42,            -- (000011.110110 | 3.84375)      => (001.01010 | 1.3125)          
    247 => 42,            -- (000011.110111 | 3.859375)     => (001.01010 | 1.3125)          
    248 => 42,            -- (000011.111000 | 3.875)        => (001.01010 | 1.3125)          
    249 => 42,            -- (000011.111001 | 3.890625)     => (001.01010 | 1.3125)          
    250 => 42,            -- (000011.111010 | 3.90625)      => (001.01010 | 1.3125)          
    251 => 42,            -- (000011.111011 | 3.921875)     => (001.01010 | 1.3125)          
    252 => 42,            -- (000011.111100 | 3.9375)       => (001.01010 | 1.3125)          
    253 => 42,            -- (000011.111101 | 3.953125)     => (001.01010 | 1.3125)          
    254 => 42,            -- (000011.111110 | 3.96875)      => (001.01010 | 1.3125)          
    255 => 42,            -- (000011.111111 | 3.984375)     => (001.01010 | 1.3125)          
    256 => 42,            -- (000100.000000 | 4.0)          => (001.01010 | 1.3125)          
    257 => 42,            -- (000100.000001 | 4.015625)     => (001.01010 | 1.3125)          
    258 => 42,            -- (000100.000010 | 4.03125)      => (001.01010 | 1.3125)          
    259 => 42,            -- (000100.000011 | 4.046875)     => (001.01010 | 1.3125)          
    260 => 42,            -- (000100.000100 | 4.0625)       => (001.01010 | 1.3125)          
    261 => 42,            -- (000100.000101 | 4.078125)     => (001.01010 | 1.3125)          
    262 => 42,            -- (000100.000110 | 4.09375)      => (001.01010 | 1.3125)          
    263 => 42,            -- (000100.000111 | 4.109375)     => (001.01010 | 1.3125)          
    264 => 42,            -- (000100.001000 | 4.125)        => (001.01010 | 1.3125)          
    265 => 42,            -- (000100.001001 | 4.140625)     => (001.01010 | 1.3125)          
    266 => 42,            -- (000100.001010 | 4.15625)      => (001.01010 | 1.3125)          
    267 => 42,            -- (000100.001011 | 4.171875)     => (001.01010 | 1.3125)          
    268 => 42,            -- (000100.001100 | 4.1875)       => (001.01010 | 1.3125)          
    269 => 42,            -- (000100.001101 | 4.203125)     => (001.01010 | 1.3125)          
    270 => 42,            -- (000100.001110 | 4.21875)      => (001.01010 | 1.3125)          
    271 => 42,            -- (000100.001111 | 4.234375)     => (001.01010 | 1.3125)          
    272 => 42,            -- (000100.010000 | 4.25)         => (001.01010 | 1.3125)          
    273 => 42,            -- (000100.010001 | 4.265625)     => (001.01010 | 1.3125)          
    274 => 42,            -- (000100.010010 | 4.28125)      => (001.01010 | 1.3125)          
    275 => 42,            -- (000100.010011 | 4.296875)     => (001.01010 | 1.3125)          
    276 => 42,            -- (000100.010100 | 4.3125)       => (001.01010 | 1.3125)          
    277 => 42,            -- (000100.010101 | 4.328125)     => (001.01010 | 1.3125)          
    278 => 43,            -- (000100.010110 | 4.34375)      => (001.01011 | 1.34375)         
    279 => 43,            -- (000100.010111 | 4.359375)     => (001.01011 | 1.34375)         
    280 => 43,            -- (000100.011000 | 4.375)        => (001.01011 | 1.34375)         
    281 => 43,            -- (000100.011001 | 4.390625)     => (001.01011 | 1.34375)         
    282 => 43,            -- (000100.011010 | 4.40625)      => (001.01011 | 1.34375)         
    283 => 43,            -- (000100.011011 | 4.421875)     => (001.01011 | 1.34375)         
    284 => 43,            -- (000100.011100 | 4.4375)       => (001.01011 | 1.34375)         
    285 => 43,            -- (000100.011101 | 4.453125)     => (001.01011 | 1.34375)         
    286 => 43,            -- (000100.011110 | 4.46875)      => (001.01011 | 1.34375)         
    287 => 43,            -- (000100.011111 | 4.484375)     => (001.01011 | 1.34375)         
    288 => 43,            -- (000100.100000 | 4.5)          => (001.01011 | 1.34375)         
    289 => 43,            -- (000100.100001 | 4.515625)     => (001.01011 | 1.34375)         
    290 => 43,            -- (000100.100010 | 4.53125)      => (001.01011 | 1.34375)         
    291 => 43,            -- (000100.100011 | 4.546875)     => (001.01011 | 1.34375)         
    292 => 43,            -- (000100.100100 | 4.5625)       => (001.01011 | 1.34375)         
    293 => 43,            -- (000100.100101 | 4.578125)     => (001.01011 | 1.34375)         
    294 => 43,            -- (000100.100110 | 4.59375)      => (001.01011 | 1.34375)         
    295 => 43,            -- (000100.100111 | 4.609375)     => (001.01011 | 1.34375)         
    296 => 43,            -- (000100.101000 | 4.625)        => (001.01011 | 1.34375)         
    297 => 43,            -- (000100.101001 | 4.640625)     => (001.01011 | 1.34375)         
    298 => 43,            -- (000100.101010 | 4.65625)      => (001.01011 | 1.34375)         
    299 => 43,            -- (000100.101011 | 4.671875)     => (001.01011 | 1.34375)         
    300 => 43,            -- (000100.101100 | 4.6875)       => (001.01011 | 1.34375)         
    301 => 43,            -- (000100.101101 | 4.703125)     => (001.01011 | 1.34375)         
    302 => 43,            -- (000100.101110 | 4.71875)      => (001.01011 | 1.34375)         
    303 => 43,            -- (000100.101111 | 4.734375)     => (001.01011 | 1.34375)         
    304 => 43,            -- (000100.110000 | 4.75)         => (001.01011 | 1.34375)         
    305 => 43,            -- (000100.110001 | 4.765625)     => (001.01011 | 1.34375)         
    306 => 43,            -- (000100.110010 | 4.78125)      => (001.01011 | 1.34375)         
    307 => 43,            -- (000100.110011 | 4.796875)     => (001.01011 | 1.34375)         
    308 => 43,            -- (000100.110100 | 4.8125)       => (001.01011 | 1.34375)         
    309 => 43,            -- (000100.110101 | 4.828125)     => (001.01011 | 1.34375)         
    310 => 43,            -- (000100.110110 | 4.84375)      => (001.01011 | 1.34375)         
    311 => 43,            -- (000100.110111 | 4.859375)     => (001.01011 | 1.34375)         
    312 => 43,            -- (000100.111000 | 4.875)        => (001.01011 | 1.34375)         
    313 => 43,            -- (000100.111001 | 4.890625)     => (001.01011 | 1.34375)         
    314 => 43,            -- (000100.111010 | 4.90625)      => (001.01011 | 1.34375)         
    315 => 43,            -- (000100.111011 | 4.921875)     => (001.01011 | 1.34375)         
    316 => 43,            -- (000100.111100 | 4.9375)       => (001.01011 | 1.34375)         
    317 => 43,            -- (000100.111101 | 4.953125)     => (001.01011 | 1.34375)         
    318 => 43,            -- (000100.111110 | 4.96875)      => (001.01011 | 1.34375)         
    319 => 43,            -- (000100.111111 | 4.984375)     => (001.01011 | 1.34375)         
    320 => 43,            -- (000101.000000 | 5.0)          => (001.01011 | 1.34375)         
    321 => 43,            -- (000101.000001 | 5.015625)     => (001.01011 | 1.34375)         
    322 => 43,            -- (000101.000010 | 5.03125)      => (001.01011 | 1.34375)         
    323 => 44,            -- (000101.000011 | 5.046875)     => (001.01100 | 1.375)           
    324 => 44,            -- (000101.000100 | 5.0625)       => (001.01100 | 1.375)           
    325 => 44,            -- (000101.000101 | 5.078125)     => (001.01100 | 1.375)           
    326 => 44,            -- (000101.000110 | 5.09375)      => (001.01100 | 1.375)           
    327 => 44,            -- (000101.000111 | 5.109375)     => (001.01100 | 1.375)           
    328 => 44,            -- (000101.001000 | 5.125)        => (001.01100 | 1.375)           
    329 => 44,            -- (000101.001001 | 5.140625)     => (001.01100 | 1.375)           
    330 => 44,            -- (000101.001010 | 5.15625)      => (001.01100 | 1.375)           
    331 => 44,            -- (000101.001011 | 5.171875)     => (001.01100 | 1.375)           
    332 => 44,            -- (000101.001100 | 5.1875)       => (001.01100 | 1.375)           
    333 => 44,            -- (000101.001101 | 5.203125)     => (001.01100 | 1.375)           
    334 => 44,            -- (000101.001110 | 5.21875)      => (001.01100 | 1.375)           
    335 => 44,            -- (000101.001111 | 5.234375)     => (001.01100 | 1.375)           
    336 => 44,            -- (000101.010000 | 5.25)         => (001.01100 | 1.375)           
    337 => 44,            -- (000101.010001 | 5.265625)     => (001.01100 | 1.375)           
    338 => 44,            -- (000101.010010 | 5.28125)      => (001.01100 | 1.375)           
    339 => 44,            -- (000101.010011 | 5.296875)     => (001.01100 | 1.375)           
    340 => 44,            -- (000101.010100 | 5.3125)       => (001.01100 | 1.375)           
    341 => 44,            -- (000101.010101 | 5.328125)     => (001.01100 | 1.375)           
    342 => 44,            -- (000101.010110 | 5.34375)      => (001.01100 | 1.375)           
    343 => 44,            -- (000101.010111 | 5.359375)     => (001.01100 | 1.375)           
    344 => 44,            -- (000101.011000 | 5.375)        => (001.01100 | 1.375)           
    345 => 44,            -- (000101.011001 | 5.390625)     => (001.01100 | 1.375)           
    346 => 44,            -- (000101.011010 | 5.40625)      => (001.01100 | 1.375)           
    347 => 44,            -- (000101.011011 | 5.421875)     => (001.01100 | 1.375)           
    348 => 44,            -- (000101.011100 | 5.4375)       => (001.01100 | 1.375)           
    349 => 44,            -- (000101.011101 | 5.453125)     => (001.01100 | 1.375)           
    350 => 44,            -- (000101.011110 | 5.46875)      => (001.01100 | 1.375)           
    351 => 44,            -- (000101.011111 | 5.484375)     => (001.01100 | 1.375)           
    352 => 44,            -- (000101.100000 | 5.5)          => (001.01100 | 1.375)           
    353 => 44,            -- (000101.100001 | 5.515625)     => (001.01100 | 1.375)           
    354 => 44,            -- (000101.100010 | 5.53125)      => (001.01100 | 1.375)           
    355 => 44,            -- (000101.100011 | 5.546875)     => (001.01100 | 1.375)           
    356 => 44,            -- (000101.100100 | 5.5625)       => (001.01100 | 1.375)           
    357 => 44,            -- (000101.100101 | 5.578125)     => (001.01100 | 1.375)           
    358 => 44,            -- (000101.100110 | 5.59375)      => (001.01100 | 1.375)           
    359 => 44,            -- (000101.100111 | 5.609375)     => (001.01100 | 1.375)           
    360 => 44,            -- (000101.101000 | 5.625)        => (001.01100 | 1.375)           
    361 => 44,            -- (000101.101001 | 5.640625)     => (001.01100 | 1.375)           
    362 => 44,            -- (000101.101010 | 5.65625)      => (001.01100 | 1.375)           
    363 => 44,            -- (000101.101011 | 5.671875)     => (001.01100 | 1.375)           
    364 => 44,            -- (000101.101100 | 5.6875)       => (001.01100 | 1.375)           
    365 => 44,            -- (000101.101101 | 5.703125)     => (001.01100 | 1.375)           
    366 => 44,            -- (000101.101110 | 5.71875)      => (001.01100 | 1.375)           
    367 => 44,            -- (000101.101111 | 5.734375)     => (001.01100 | 1.375)           
    368 => 44,            -- (000101.110000 | 5.75)         => (001.01100 | 1.375)           
    369 => 44,            -- (000101.110001 | 5.765625)     => (001.01100 | 1.375)           
    370 => 44,            -- (000101.110010 | 5.78125)      => (001.01100 | 1.375)           
    371 => 44,            -- (000101.110011 | 5.796875)     => (001.01100 | 1.375)           
    372 => 44,            -- (000101.110100 | 5.8125)       => (001.01100 | 1.375)           
    373 => 44,            -- (000101.110101 | 5.828125)     => (001.01100 | 1.375)           
    374 => 44,            -- (000101.110110 | 5.84375)      => (001.01100 | 1.375)           
    375 => 44,            -- (000101.110111 | 5.859375)     => (001.01100 | 1.375)           
    376 => 44,            -- (000101.111000 | 5.875)        => (001.01100 | 1.375)           
    377 => 44,            -- (000101.111001 | 5.890625)     => (001.01100 | 1.375)           
    378 => 44,            -- (000101.111010 | 5.90625)      => (001.01100 | 1.375)           
    379 => 44,            -- (000101.111011 | 5.921875)     => (001.01100 | 1.375)           
    380 => 44,            -- (000101.111100 | 5.9375)       => (001.01100 | 1.375)           
    381 => 44,            -- (000101.111101 | 5.953125)     => (001.01100 | 1.375)           
    382 => 44,            -- (000101.111110 | 5.96875)      => (001.01100 | 1.375)           
    383 => 44,            -- (000101.111111 | 5.984375)     => (001.01100 | 1.375)           
    384 => 44,            -- (000110.000000 | 6.0)          => (001.01100 | 1.375)           
    385 => 44,            -- (000110.000001 | 6.015625)     => (001.01100 | 1.375)           
    386 => 45,            -- (000110.000010 | 6.03125)      => (001.01101 | 1.40625)         
    387 => 45,            -- (000110.000011 | 6.046875)     => (001.01101 | 1.40625)         
    388 => 45,            -- (000110.000100 | 6.0625)       => (001.01101 | 1.40625)         
    389 => 45,            -- (000110.000101 | 6.078125)     => (001.01101 | 1.40625)         
    390 => 45,            -- (000110.000110 | 6.09375)      => (001.01101 | 1.40625)         
    391 => 45,            -- (000110.000111 | 6.109375)     => (001.01101 | 1.40625)         
    392 => 45,            -- (000110.001000 | 6.125)        => (001.01101 | 1.40625)         
    393 => 45,            -- (000110.001001 | 6.140625)     => (001.01101 | 1.40625)         
    394 => 45,            -- (000110.001010 | 6.15625)      => (001.01101 | 1.40625)         
    395 => 45,            -- (000110.001011 | 6.171875)     => (001.01101 | 1.40625)         
    396 => 45,            -- (000110.001100 | 6.1875)       => (001.01101 | 1.40625)         
    397 => 45,            -- (000110.001101 | 6.203125)     => (001.01101 | 1.40625)         
    398 => 45,            -- (000110.001110 | 6.21875)      => (001.01101 | 1.40625)         
    399 => 45,            -- (000110.001111 | 6.234375)     => (001.01101 | 1.40625)         
    400 => 45,            -- (000110.010000 | 6.25)         => (001.01101 | 1.40625)         
    401 => 45,            -- (000110.010001 | 6.265625)     => (001.01101 | 1.40625)         
    402 => 45,            -- (000110.010010 | 6.28125)      => (001.01101 | 1.40625)         
    403 => 45,            -- (000110.010011 | 6.296875)     => (001.01101 | 1.40625)         
    404 => 45,            -- (000110.010100 | 6.3125)       => (001.01101 | 1.40625)         
    405 => 45,            -- (000110.010101 | 6.328125)     => (001.01101 | 1.40625)         
    406 => 45,            -- (000110.010110 | 6.34375)      => (001.01101 | 1.40625)         
    407 => 45,            -- (000110.010111 | 6.359375)     => (001.01101 | 1.40625)         
    408 => 45,            -- (000110.011000 | 6.375)        => (001.01101 | 1.40625)         
    409 => 45,            -- (000110.011001 | 6.390625)     => (001.01101 | 1.40625)         
    410 => 45,            -- (000110.011010 | 6.40625)      => (001.01101 | 1.40625)         
    411 => 45,            -- (000110.011011 | 6.421875)     => (001.01101 | 1.40625)         
    412 => 45,            -- (000110.011100 | 6.4375)       => (001.01101 | 1.40625)         
    413 => 45,            -- (000110.011101 | 6.453125)     => (001.01101 | 1.40625)         
    414 => 45,            -- (000110.011110 | 6.46875)      => (001.01101 | 1.40625)         
    415 => 45,            -- (000110.011111 | 6.484375)     => (001.01101 | 1.40625)         
    416 => 45,            -- (000110.100000 | 6.5)          => (001.01101 | 1.40625)         
    417 => 45,            -- (000110.100001 | 6.515625)     => (001.01101 | 1.40625)         
    418 => 45,            -- (000110.100010 | 6.53125)      => (001.01101 | 1.40625)         
    419 => 45,            -- (000110.100011 | 6.546875)     => (001.01101 | 1.40625)         
    420 => 45,            -- (000110.100100 | 6.5625)       => (001.01101 | 1.40625)         
    421 => 45,            -- (000110.100101 | 6.578125)     => (001.01101 | 1.40625)         
    422 => 45,            -- (000110.100110 | 6.59375)      => (001.01101 | 1.40625)         
    423 => 45,            -- (000110.100111 | 6.609375)     => (001.01101 | 1.40625)         
    424 => 45,            -- (000110.101000 | 6.625)        => (001.01101 | 1.40625)         
    425 => 45,            -- (000110.101001 | 6.640625)     => (001.01101 | 1.40625)         
    426 => 45,            -- (000110.101010 | 6.65625)      => (001.01101 | 1.40625)         
    427 => 45,            -- (000110.101011 | 6.671875)     => (001.01101 | 1.40625)         
    428 => 45,            -- (000110.101100 | 6.6875)       => (001.01101 | 1.40625)         
    429 => 45,            -- (000110.101101 | 6.703125)     => (001.01101 | 1.40625)         
    430 => 45,            -- (000110.101110 | 6.71875)      => (001.01101 | 1.40625)         
    431 => 45,            -- (000110.101111 | 6.734375)     => (001.01101 | 1.40625)         
    432 => 45,            -- (000110.110000 | 6.75)         => (001.01101 | 1.40625)         
    433 => 45,            -- (000110.110001 | 6.765625)     => (001.01101 | 1.40625)         
    434 => 45,            -- (000110.110010 | 6.78125)      => (001.01101 | 1.40625)         
    435 => 45,            -- (000110.110011 | 6.796875)     => (001.01101 | 1.40625)         
    436 => 45,            -- (000110.110100 | 6.8125)       => (001.01101 | 1.40625)         
    437 => 45,            -- (000110.110101 | 6.828125)     => (001.01101 | 1.40625)         
    438 => 45,            -- (000110.110110 | 6.84375)      => (001.01101 | 1.40625)         
    439 => 45,            -- (000110.110111 | 6.859375)     => (001.01101 | 1.40625)         
    440 => 45,            -- (000110.111000 | 6.875)        => (001.01101 | 1.40625)         
    441 => 45,            -- (000110.111001 | 6.890625)     => (001.01101 | 1.40625)         
    442 => 45,            -- (000110.111010 | 6.90625)      => (001.01101 | 1.40625)         
    443 => 45,            -- (000110.111011 | 6.921875)     => (001.01101 | 1.40625)         
    444 => 45,            -- (000110.111100 | 6.9375)       => (001.01101 | 1.40625)         
    445 => 45,            -- (000110.111101 | 6.953125)     => (001.01101 | 1.40625)         
    446 => 45,            -- (000110.111110 | 6.96875)      => (001.01101 | 1.40625)         
    447 => 45,            -- (000110.111111 | 6.984375)     => (001.01101 | 1.40625)         
    448 => 45,            -- (000111.000000 | 7.0)          => (001.01101 | 1.40625)         
    449 => 45,            -- (000111.000001 | 7.015625)     => (001.01101 | 1.40625)         
    450 => 45,            -- (000111.000010 | 7.03125)      => (001.01101 | 1.40625)         
    451 => 45,            -- (000111.000011 | 7.046875)     => (001.01101 | 1.40625)         
    452 => 45,            -- (000111.000100 | 7.0625)       => (001.01101 | 1.40625)         
    453 => 45,            -- (000111.000101 | 7.078125)     => (001.01101 | 1.40625)         
    454 => 45,            -- (000111.000110 | 7.09375)      => (001.01101 | 1.40625)         
    455 => 45,            -- (000111.000111 | 7.109375)     => (001.01101 | 1.40625)         
    456 => 45,            -- (000111.001000 | 7.125)        => (001.01101 | 1.40625)         
    457 => 45,            -- (000111.001001 | 7.140625)     => (001.01101 | 1.40625)         
    458 => 45,            -- (000111.001010 | 7.15625)      => (001.01101 | 1.40625)         
    459 => 45,            -- (000111.001011 | 7.171875)     => (001.01101 | 1.40625)         
    460 => 45,            -- (000111.001100 | 7.1875)       => (001.01101 | 1.40625)         
    461 => 45,            -- (000111.001101 | 7.203125)     => (001.01101 | 1.40625)         
    462 => 45,            -- (000111.001110 | 7.21875)      => (001.01101 | 1.40625)         
    463 => 45,            -- (000111.001111 | 7.234375)     => (001.01101 | 1.40625)         
    464 => 45,            -- (000111.010000 | 7.25)         => (001.01101 | 1.40625)         
    465 => 45,            -- (000111.010001 | 7.265625)     => (001.01101 | 1.40625)         
    466 => 45,            -- (000111.010010 | 7.28125)      => (001.01101 | 1.40625)         
    467 => 45,            -- (000111.010011 | 7.296875)     => (001.01101 | 1.40625)         
    468 => 45,            -- (000111.010100 | 7.3125)       => (001.01101 | 1.40625)         
    469 => 45,            -- (000111.010101 | 7.328125)     => (001.01101 | 1.40625)         
    470 => 45,            -- (000111.010110 | 7.34375)      => (001.01101 | 1.40625)         
    471 => 45,            -- (000111.010111 | 7.359375)     => (001.01101 | 1.40625)         
    472 => 45,            -- (000111.011000 | 7.375)        => (001.01101 | 1.40625)         
    473 => 45,            -- (000111.011001 | 7.390625)     => (001.01101 | 1.40625)         
    474 => 45,            -- (000111.011010 | 7.40625)      => (001.01101 | 1.40625)         
    475 => 45,            -- (000111.011011 | 7.421875)     => (001.01101 | 1.40625)         
    476 => 45,            -- (000111.011100 | 7.4375)       => (001.01101 | 1.40625)         
    477 => 45,            -- (000111.011101 | 7.453125)     => (001.01101 | 1.40625)         
    478 => 46,            -- (000111.011110 | 7.46875)      => (001.01110 | 1.4375)          
    479 => 46,            -- (000111.011111 | 7.484375)     => (001.01110 | 1.4375)          
    480 => 46,            -- (000111.100000 | 7.5)          => (001.01110 | 1.4375)          
    481 => 46,            -- (000111.100001 | 7.515625)     => (001.01110 | 1.4375)          
    482 => 46,            -- (000111.100010 | 7.53125)      => (001.01110 | 1.4375)          
    483 => 46,            -- (000111.100011 | 7.546875)     => (001.01110 | 1.4375)          
    484 => 46,            -- (000111.100100 | 7.5625)       => (001.01110 | 1.4375)          
    485 => 46,            -- (000111.100101 | 7.578125)     => (001.01110 | 1.4375)          
    486 => 46,            -- (000111.100110 | 7.59375)      => (001.01110 | 1.4375)          
    487 => 46,            -- (000111.100111 | 7.609375)     => (001.01110 | 1.4375)          
    488 => 46,            -- (000111.101000 | 7.625)        => (001.01110 | 1.4375)          
    489 => 46,            -- (000111.101001 | 7.640625)     => (001.01110 | 1.4375)          
    490 => 46,            -- (000111.101010 | 7.65625)      => (001.01110 | 1.4375)          
    491 => 46,            -- (000111.101011 | 7.671875)     => (001.01110 | 1.4375)          
    492 => 46,            -- (000111.101100 | 7.6875)       => (001.01110 | 1.4375)          
    493 => 46,            -- (000111.101101 | 7.703125)     => (001.01110 | 1.4375)          
    494 => 46,            -- (000111.101110 | 7.71875)      => (001.01110 | 1.4375)          
    495 => 46,            -- (000111.101111 | 7.734375)     => (001.01110 | 1.4375)          
    496 => 46,            -- (000111.110000 | 7.75)         => (001.01110 | 1.4375)          
    497 => 46,            -- (000111.110001 | 7.765625)     => (001.01110 | 1.4375)          
    498 => 46,            -- (000111.110010 | 7.78125)      => (001.01110 | 1.4375)          
    499 => 46,            -- (000111.110011 | 7.796875)     => (001.01110 | 1.4375)          
    500 => 46,            -- (000111.110100 | 7.8125)       => (001.01110 | 1.4375)          
    501 => 46,            -- (000111.110101 | 7.828125)     => (001.01110 | 1.4375)          
    502 => 46,            -- (000111.110110 | 7.84375)      => (001.01110 | 1.4375)          
    503 => 46,            -- (000111.110111 | 7.859375)     => (001.01110 | 1.4375)          
    504 => 46,            -- (000111.111000 | 7.875)        => (001.01110 | 1.4375)          
    505 => 46,            -- (000111.111001 | 7.890625)     => (001.01110 | 1.4375)          
    506 => 46,            -- (000111.111010 | 7.90625)      => (001.01110 | 1.4375)          
    507 => 46,            -- (000111.111011 | 7.921875)     => (001.01110 | 1.4375)          
    508 => 46,            -- (000111.111100 | 7.9375)       => (001.01110 | 1.4375)          
    509 => 46,            -- (000111.111101 | 7.953125)     => (001.01110 | 1.4375)          
    510 => 46,            -- (000111.111110 | 7.96875)      => (001.01110 | 1.4375)          
    511 => 46,            -- (000111.111111 | 7.984375)     => (001.01110 | 1.4375)          
    512 => 46,            -- (001000.000000 | 8.0)          => (001.01110 | 1.4375)          
    513 => 46,            -- (001000.000001 | 8.015625)     => (001.01110 | 1.4375)          
    514 => 46,            -- (001000.000010 | 8.03125)      => (001.01110 | 1.4375)          
    515 => 46,            -- (001000.000011 | 8.046875)     => (001.01110 | 1.4375)          
    516 => 46,            -- (001000.000100 | 8.0625)       => (001.01110 | 1.4375)          
    517 => 46,            -- (001000.000101 | 8.078125)     => (001.01110 | 1.4375)          
    518 => 46,            -- (001000.000110 | 8.09375)      => (001.01110 | 1.4375)          
    519 => 46,            -- (001000.000111 | 8.109375)     => (001.01110 | 1.4375)          
    520 => 46,            -- (001000.001000 | 8.125)        => (001.01110 | 1.4375)          
    521 => 46,            -- (001000.001001 | 8.140625)     => (001.01110 | 1.4375)          
    522 => 46,            -- (001000.001010 | 8.15625)      => (001.01110 | 1.4375)          
    523 => 46,            -- (001000.001011 | 8.171875)     => (001.01110 | 1.4375)          
    524 => 46,            -- (001000.001100 | 8.1875)       => (001.01110 | 1.4375)          
    525 => 46,            -- (001000.001101 | 8.203125)     => (001.01110 | 1.4375)          
    526 => 46,            -- (001000.001110 | 8.21875)      => (001.01110 | 1.4375)          
    527 => 46,            -- (001000.001111 | 8.234375)     => (001.01110 | 1.4375)          
    528 => 46,            -- (001000.010000 | 8.25)         => (001.01110 | 1.4375)          
    529 => 46,            -- (001000.010001 | 8.265625)     => (001.01110 | 1.4375)          
    530 => 46,            -- (001000.010010 | 8.28125)      => (001.01110 | 1.4375)          
    531 => 46,            -- (001000.010011 | 8.296875)     => (001.01110 | 1.4375)          
    532 => 46,            -- (001000.010100 | 8.3125)       => (001.01110 | 1.4375)          
    533 => 46,            -- (001000.010101 | 8.328125)     => (001.01110 | 1.4375)          
    534 => 46,            -- (001000.010110 | 8.34375)      => (001.01110 | 1.4375)          
    535 => 46,            -- (001000.010111 | 8.359375)     => (001.01110 | 1.4375)          
    536 => 46,            -- (001000.011000 | 8.375)        => (001.01110 | 1.4375)          
    537 => 46,            -- (001000.011001 | 8.390625)     => (001.01110 | 1.4375)          
    538 => 46,            -- (001000.011010 | 8.40625)      => (001.01110 | 1.4375)          
    539 => 46,            -- (001000.011011 | 8.421875)     => (001.01110 | 1.4375)          
    540 => 46,            -- (001000.011100 | 8.4375)       => (001.01110 | 1.4375)          
    541 => 46,            -- (001000.011101 | 8.453125)     => (001.01110 | 1.4375)          
    542 => 46,            -- (001000.011110 | 8.46875)      => (001.01110 | 1.4375)          
    543 => 46,            -- (001000.011111 | 8.484375)     => (001.01110 | 1.4375)          
    544 => 46,            -- (001000.100000 | 8.5)          => (001.01110 | 1.4375)          
    545 => 46,            -- (001000.100001 | 8.515625)     => (001.01110 | 1.4375)          
    546 => 46,            -- (001000.100010 | 8.53125)      => (001.01110 | 1.4375)          
    547 => 46,            -- (001000.100011 | 8.546875)     => (001.01110 | 1.4375)          
    548 => 46,            -- (001000.100100 | 8.5625)       => (001.01110 | 1.4375)          
    549 => 46,            -- (001000.100101 | 8.578125)     => (001.01110 | 1.4375)          
    550 => 46,            -- (001000.100110 | 8.59375)      => (001.01110 | 1.4375)          
    551 => 46,            -- (001000.100111 | 8.609375)     => (001.01110 | 1.4375)          
    552 => 46,            -- (001000.101000 | 8.625)        => (001.01110 | 1.4375)          
    553 => 46,            -- (001000.101001 | 8.640625)     => (001.01110 | 1.4375)          
    554 => 46,            -- (001000.101010 | 8.65625)      => (001.01110 | 1.4375)          
    555 => 46,            -- (001000.101011 | 8.671875)     => (001.01110 | 1.4375)          
    556 => 46,            -- (001000.101100 | 8.6875)       => (001.01110 | 1.4375)          
    557 => 46,            -- (001000.101101 | 8.703125)     => (001.01110 | 1.4375)          
    558 => 46,            -- (001000.101110 | 8.71875)      => (001.01110 | 1.4375)          
    559 => 46,            -- (001000.101111 | 8.734375)     => (001.01110 | 1.4375)          
    560 => 46,            -- (001000.110000 | 8.75)         => (001.01110 | 1.4375)          
    561 => 46,            -- (001000.110001 | 8.765625)     => (001.01110 | 1.4375)          
    562 => 46,            -- (001000.110010 | 8.78125)      => (001.01110 | 1.4375)          
    563 => 46,            -- (001000.110011 | 8.796875)     => (001.01110 | 1.4375)          
    564 => 46,            -- (001000.110100 | 8.8125)       => (001.01110 | 1.4375)          
    565 => 46,            -- (001000.110101 | 8.828125)     => (001.01110 | 1.4375)          
    566 => 46,            -- (001000.110110 | 8.84375)      => (001.01110 | 1.4375)          
    567 => 46,            -- (001000.110111 | 8.859375)     => (001.01110 | 1.4375)          
    568 => 46,            -- (001000.111000 | 8.875)        => (001.01110 | 1.4375)          
    569 => 46,            -- (001000.111001 | 8.890625)     => (001.01110 | 1.4375)          
    570 => 46,            -- (001000.111010 | 8.90625)      => (001.01110 | 1.4375)          
    571 => 46,            -- (001000.111011 | 8.921875)     => (001.01110 | 1.4375)          
    572 => 46,            -- (001000.111100 | 8.9375)       => (001.01110 | 1.4375)          
    573 => 46,            -- (001000.111101 | 8.953125)     => (001.01110 | 1.4375)          
    574 => 46,            -- (001000.111110 | 8.96875)      => (001.01110 | 1.4375)          
    575 => 46,            -- (001000.111111 | 8.984375)     => (001.01110 | 1.4375)          
    576 => 46,            -- (001001.000000 | 9.0)          => (001.01110 | 1.4375)          
    577 => 46,            -- (001001.000001 | 9.015625)     => (001.01110 | 1.4375)          
    578 => 46,            -- (001001.000010 | 9.03125)      => (001.01110 | 1.4375)          
    579 => 46,            -- (001001.000011 | 9.046875)     => (001.01110 | 1.4375)          
    580 => 46,            -- (001001.000100 | 9.0625)       => (001.01110 | 1.4375)          
    581 => 46,            -- (001001.000101 | 9.078125)     => (001.01110 | 1.4375)          
    582 => 46,            -- (001001.000110 | 9.09375)      => (001.01110 | 1.4375)          
    583 => 46,            -- (001001.000111 | 9.109375)     => (001.01110 | 1.4375)          
    584 => 46,            -- (001001.001000 | 9.125)        => (001.01110 | 1.4375)          
    585 => 46,            -- (001001.001001 | 9.140625)     => (001.01110 | 1.4375)          
    586 => 46,            -- (001001.001010 | 9.15625)      => (001.01110 | 1.4375)          
    587 => 46,            -- (001001.001011 | 9.171875)     => (001.01110 | 1.4375)          
    588 => 46,            -- (001001.001100 | 9.1875)       => (001.01110 | 1.4375)          
    589 => 46,            -- (001001.001101 | 9.203125)     => (001.01110 | 1.4375)          
    590 => 46,            -- (001001.001110 | 9.21875)      => (001.01110 | 1.4375)          
    591 => 46,            -- (001001.001111 | 9.234375)     => (001.01110 | 1.4375)          
    592 => 46,            -- (001001.010000 | 9.25)         => (001.01110 | 1.4375)          
    593 => 46,            -- (001001.010001 | 9.265625)     => (001.01110 | 1.4375)          
    594 => 46,            -- (001001.010010 | 9.28125)      => (001.01110 | 1.4375)          
    595 => 46,            -- (001001.010011 | 9.296875)     => (001.01110 | 1.4375)          
    596 => 46,            -- (001001.010100 | 9.3125)       => (001.01110 | 1.4375)          
    597 => 46,            -- (001001.010101 | 9.328125)     => (001.01110 | 1.4375)          
    598 => 46,            -- (001001.010110 | 9.34375)      => (001.01110 | 1.4375)          
    599 => 46,            -- (001001.010111 | 9.359375)     => (001.01110 | 1.4375)          
    600 => 46,            -- (001001.011000 | 9.375)        => (001.01110 | 1.4375)          
    601 => 46,            -- (001001.011001 | 9.390625)     => (001.01110 | 1.4375)          
    602 => 46,            -- (001001.011010 | 9.40625)      => (001.01110 | 1.4375)          
    603 => 46,            -- (001001.011011 | 9.421875)     => (001.01110 | 1.4375)          
    604 => 46,            -- (001001.011100 | 9.4375)       => (001.01110 | 1.4375)          
    605 => 46,            -- (001001.011101 | 9.453125)     => (001.01110 | 1.4375)          
    606 => 46,            -- (001001.011110 | 9.46875)      => (001.01110 | 1.4375)          
    607 => 46,            -- (001001.011111 | 9.484375)     => (001.01110 | 1.4375)          
    608 => 46,            -- (001001.100000 | 9.5)          => (001.01110 | 1.4375)          
    609 => 46,            -- (001001.100001 | 9.515625)     => (001.01110 | 1.4375)          
    610 => 46,            -- (001001.100010 | 9.53125)      => (001.01110 | 1.4375)          
    611 => 46,            -- (001001.100011 | 9.546875)     => (001.01110 | 1.4375)          
    612 => 46,            -- (001001.100100 | 9.5625)       => (001.01110 | 1.4375)          
    613 => 46,            -- (001001.100101 | 9.578125)     => (001.01110 | 1.4375)          
    614 => 46,            -- (001001.100110 | 9.59375)      => (001.01110 | 1.4375)          
    615 => 46,            -- (001001.100111 | 9.609375)     => (001.01110 | 1.4375)          
    616 => 46,            -- (001001.101000 | 9.625)        => (001.01110 | 1.4375)          
    617 => 46,            -- (001001.101001 | 9.640625)     => (001.01110 | 1.4375)          
    618 => 46,            -- (001001.101010 | 9.65625)      => (001.01110 | 1.4375)          
    619 => 46,            -- (001001.101011 | 9.671875)     => (001.01110 | 1.4375)          
    620 => 46,            -- (001001.101100 | 9.6875)       => (001.01110 | 1.4375)          
    621 => 46,            -- (001001.101101 | 9.703125)     => (001.01110 | 1.4375)          
    622 => 46,            -- (001001.101110 | 9.71875)      => (001.01110 | 1.4375)          
    623 => 46,            -- (001001.101111 | 9.734375)     => (001.01110 | 1.4375)          
    624 => 46,            -- (001001.110000 | 9.75)         => (001.01110 | 1.4375)          
    625 => 47,            -- (001001.110001 | 9.765625)     => (001.01111 | 1.46875)         
    626 => 47,            -- (001001.110010 | 9.78125)      => (001.01111 | 1.46875)         
    627 => 47,            -- (001001.110011 | 9.796875)     => (001.01111 | 1.46875)         
    628 => 47,            -- (001001.110100 | 9.8125)       => (001.01111 | 1.46875)         
    629 => 47,            -- (001001.110101 | 9.828125)     => (001.01111 | 1.46875)         
    630 => 47,            -- (001001.110110 | 9.84375)      => (001.01111 | 1.46875)         
    631 => 47,            -- (001001.110111 | 9.859375)     => (001.01111 | 1.46875)         
    632 => 47,            -- (001001.111000 | 9.875)        => (001.01111 | 1.46875)         
    633 => 47,            -- (001001.111001 | 9.890625)     => (001.01111 | 1.46875)         
    634 => 47,            -- (001001.111010 | 9.90625)      => (001.01111 | 1.46875)         
    635 => 47,            -- (001001.111011 | 9.921875)     => (001.01111 | 1.46875)         
    636 => 47,            -- (001001.111100 | 9.9375)       => (001.01111 | 1.46875)         
    637 => 47,            -- (001001.111101 | 9.953125)     => (001.01111 | 1.46875)         
    638 => 47,            -- (001001.111110 | 9.96875)      => (001.01111 | 1.46875)         
    639 => 47,            -- (001001.111111 | 9.984375)     => (001.01111 | 1.46875)         
    640 => 47,            -- (001010.000000 | 10.0)         => (001.01111 | 1.46875)         
    641 => 47,            -- (001010.000001 | 10.015625)    => (001.01111 | 1.46875)         
    642 => 47,            -- (001010.000010 | 10.03125)     => (001.01111 | 1.46875)         
    643 => 47,            -- (001010.000011 | 10.046875)    => (001.01111 | 1.46875)         
    644 => 47,            -- (001010.000100 | 10.0625)      => (001.01111 | 1.46875)         
    645 => 47,            -- (001010.000101 | 10.078125)    => (001.01111 | 1.46875)         
    646 => 47,            -- (001010.000110 | 10.09375)     => (001.01111 | 1.46875)         
    647 => 47,            -- (001010.000111 | 10.109375)    => (001.01111 | 1.46875)         
    648 => 47,            -- (001010.001000 | 10.125)       => (001.01111 | 1.46875)         
    649 => 47,            -- (001010.001001 | 10.140625)    => (001.01111 | 1.46875)         
    650 => 47,            -- (001010.001010 | 10.15625)     => (001.01111 | 1.46875)         
    651 => 47,            -- (001010.001011 | 10.171875)    => (001.01111 | 1.46875)         
    652 => 47,            -- (001010.001100 | 10.1875)      => (001.01111 | 1.46875)         
    653 => 47,            -- (001010.001101 | 10.203125)    => (001.01111 | 1.46875)         
    654 => 47,            -- (001010.001110 | 10.21875)     => (001.01111 | 1.46875)         
    655 => 47,            -- (001010.001111 | 10.234375)    => (001.01111 | 1.46875)         
    656 => 47,            -- (001010.010000 | 10.25)        => (001.01111 | 1.46875)         
    657 => 47,            -- (001010.010001 | 10.265625)    => (001.01111 | 1.46875)         
    658 => 47,            -- (001010.010010 | 10.28125)     => (001.01111 | 1.46875)         
    659 => 47,            -- (001010.010011 | 10.296875)    => (001.01111 | 1.46875)         
    660 => 47,            -- (001010.010100 | 10.3125)      => (001.01111 | 1.46875)         
    661 => 47,            -- (001010.010101 | 10.328125)    => (001.01111 | 1.46875)         
    662 => 47,            -- (001010.010110 | 10.34375)     => (001.01111 | 1.46875)         
    663 => 47,            -- (001010.010111 | 10.359375)    => (001.01111 | 1.46875)         
    664 => 47,            -- (001010.011000 | 10.375)       => (001.01111 | 1.46875)         
    665 => 47,            -- (001010.011001 | 10.390625)    => (001.01111 | 1.46875)         
    666 => 47,            -- (001010.011010 | 10.40625)     => (001.01111 | 1.46875)         
    667 => 47,            -- (001010.011011 | 10.421875)    => (001.01111 | 1.46875)         
    668 => 47,            -- (001010.011100 | 10.4375)      => (001.01111 | 1.46875)         
    669 => 47,            -- (001010.011101 | 10.453125)    => (001.01111 | 1.46875)         
    670 => 47,            -- (001010.011110 | 10.46875)     => (001.01111 | 1.46875)         
    671 => 47,            -- (001010.011111 | 10.484375)    => (001.01111 | 1.46875)         
    672 => 47,            -- (001010.100000 | 10.5)         => (001.01111 | 1.46875)         
    673 => 47,            -- (001010.100001 | 10.515625)    => (001.01111 | 1.46875)         
    674 => 47,            -- (001010.100010 | 10.53125)     => (001.01111 | 1.46875)         
    675 => 47,            -- (001010.100011 | 10.546875)    => (001.01111 | 1.46875)         
    676 => 47,            -- (001010.100100 | 10.5625)      => (001.01111 | 1.46875)         
    677 => 47,            -- (001010.100101 | 10.578125)    => (001.01111 | 1.46875)         
    678 => 47,            -- (001010.100110 | 10.59375)     => (001.01111 | 1.46875)         
    679 => 47,            -- (001010.100111 | 10.609375)    => (001.01111 | 1.46875)         
    680 => 47,            -- (001010.101000 | 10.625)       => (001.01111 | 1.46875)         
    681 => 47,            -- (001010.101001 | 10.640625)    => (001.01111 | 1.46875)         
    682 => 47,            -- (001010.101010 | 10.65625)     => (001.01111 | 1.46875)         
    683 => 47,            -- (001010.101011 | 10.671875)    => (001.01111 | 1.46875)         
    684 => 47,            -- (001010.101100 | 10.6875)      => (001.01111 | 1.46875)         
    685 => 47,            -- (001010.101101 | 10.703125)    => (001.01111 | 1.46875)         
    686 => 47,            -- (001010.101110 | 10.71875)     => (001.01111 | 1.46875)         
    687 => 47,            -- (001010.101111 | 10.734375)    => (001.01111 | 1.46875)         
    688 => 47,            -- (001010.110000 | 10.75)        => (001.01111 | 1.46875)         
    689 => 47,            -- (001010.110001 | 10.765625)    => (001.01111 | 1.46875)         
    690 => 47,            -- (001010.110010 | 10.78125)     => (001.01111 | 1.46875)         
    691 => 47,            -- (001010.110011 | 10.796875)    => (001.01111 | 1.46875)         
    692 => 47,            -- (001010.110100 | 10.8125)      => (001.01111 | 1.46875)         
    693 => 47,            -- (001010.110101 | 10.828125)    => (001.01111 | 1.46875)         
    694 => 47,            -- (001010.110110 | 10.84375)     => (001.01111 | 1.46875)         
    695 => 47,            -- (001010.110111 | 10.859375)    => (001.01111 | 1.46875)         
    696 => 47,            -- (001010.111000 | 10.875)       => (001.01111 | 1.46875)         
    697 => 47,            -- (001010.111001 | 10.890625)    => (001.01111 | 1.46875)         
    698 => 47,            -- (001010.111010 | 10.90625)     => (001.01111 | 1.46875)         
    699 => 47,            -- (001010.111011 | 10.921875)    => (001.01111 | 1.46875)         
    700 => 47,            -- (001010.111100 | 10.9375)      => (001.01111 | 1.46875)         
    701 => 47,            -- (001010.111101 | 10.953125)    => (001.01111 | 1.46875)         
    702 => 47,            -- (001010.111110 | 10.96875)     => (001.01111 | 1.46875)         
    703 => 47,            -- (001010.111111 | 10.984375)    => (001.01111 | 1.46875)         
    704 => 47,            -- (001011.000000 | 11.0)         => (001.01111 | 1.46875)         
    705 => 47,            -- (001011.000001 | 11.015625)    => (001.01111 | 1.46875)         
    706 => 47,            -- (001011.000010 | 11.03125)     => (001.01111 | 1.46875)         
    707 => 47,            -- (001011.000011 | 11.046875)    => (001.01111 | 1.46875)         
    708 => 47,            -- (001011.000100 | 11.0625)      => (001.01111 | 1.46875)         
    709 => 47,            -- (001011.000101 | 11.078125)    => (001.01111 | 1.46875)         
    710 => 47,            -- (001011.000110 | 11.09375)     => (001.01111 | 1.46875)         
    711 => 47,            -- (001011.000111 | 11.109375)    => (001.01111 | 1.46875)         
    712 => 47,            -- (001011.001000 | 11.125)       => (001.01111 | 1.46875)         
    713 => 47,            -- (001011.001001 | 11.140625)    => (001.01111 | 1.46875)         
    714 => 47,            -- (001011.001010 | 11.15625)     => (001.01111 | 1.46875)         
    715 => 47,            -- (001011.001011 | 11.171875)    => (001.01111 | 1.46875)         
    716 => 47,            -- (001011.001100 | 11.1875)      => (001.01111 | 1.46875)         
    717 => 47,            -- (001011.001101 | 11.203125)    => (001.01111 | 1.46875)         
    718 => 47,            -- (001011.001110 | 11.21875)     => (001.01111 | 1.46875)         
    719 => 47,            -- (001011.001111 | 11.234375)    => (001.01111 | 1.46875)         
    720 => 47,            -- (001011.010000 | 11.25)        => (001.01111 | 1.46875)         
    721 => 47,            -- (001011.010001 | 11.265625)    => (001.01111 | 1.46875)         
    722 => 47,            -- (001011.010010 | 11.28125)     => (001.01111 | 1.46875)         
    723 => 47,            -- (001011.010011 | 11.296875)    => (001.01111 | 1.46875)         
    724 => 47,            -- (001011.010100 | 11.3125)      => (001.01111 | 1.46875)         
    725 => 47,            -- (001011.010101 | 11.328125)    => (001.01111 | 1.46875)         
    726 => 47,            -- (001011.010110 | 11.34375)     => (001.01111 | 1.46875)         
    727 => 47,            -- (001011.010111 | 11.359375)    => (001.01111 | 1.46875)         
    728 => 47,            -- (001011.011000 | 11.375)       => (001.01111 | 1.46875)         
    729 => 47,            -- (001011.011001 | 11.390625)    => (001.01111 | 1.46875)         
    730 => 47,            -- (001011.011010 | 11.40625)     => (001.01111 | 1.46875)         
    731 => 47,            -- (001011.011011 | 11.421875)    => (001.01111 | 1.46875)         
    732 => 47,            -- (001011.011100 | 11.4375)      => (001.01111 | 1.46875)         
    733 => 47,            -- (001011.011101 | 11.453125)    => (001.01111 | 1.46875)         
    734 => 47,            -- (001011.011110 | 11.46875)     => (001.01111 | 1.46875)         
    735 => 47,            -- (001011.011111 | 11.484375)    => (001.01111 | 1.46875)         
    736 => 47,            -- (001011.100000 | 11.5)         => (001.01111 | 1.46875)         
    737 => 47,            -- (001011.100001 | 11.515625)    => (001.01111 | 1.46875)         
    738 => 47,            -- (001011.100010 | 11.53125)     => (001.01111 | 1.46875)         
    739 => 47,            -- (001011.100011 | 11.546875)    => (001.01111 | 1.46875)         
    740 => 47,            -- (001011.100100 | 11.5625)      => (001.01111 | 1.46875)         
    741 => 47,            -- (001011.100101 | 11.578125)    => (001.01111 | 1.46875)         
    742 => 47,            -- (001011.100110 | 11.59375)     => (001.01111 | 1.46875)         
    743 => 47,            -- (001011.100111 | 11.609375)    => (001.01111 | 1.46875)         
    744 => 47,            -- (001011.101000 | 11.625)       => (001.01111 | 1.46875)         
    745 => 47,            -- (001011.101001 | 11.640625)    => (001.01111 | 1.46875)         
    746 => 47,            -- (001011.101010 | 11.65625)     => (001.01111 | 1.46875)         
    747 => 47,            -- (001011.101011 | 11.671875)    => (001.01111 | 1.46875)         
    748 => 47,            -- (001011.101100 | 11.6875)      => (001.01111 | 1.46875)         
    749 => 47,            -- (001011.101101 | 11.703125)    => (001.01111 | 1.46875)         
    750 => 47,            -- (001011.101110 | 11.71875)     => (001.01111 | 1.46875)         
    751 => 47,            -- (001011.101111 | 11.734375)    => (001.01111 | 1.46875)         
    752 => 47,            -- (001011.110000 | 11.75)        => (001.01111 | 1.46875)         
    753 => 47,            -- (001011.110001 | 11.765625)    => (001.01111 | 1.46875)         
    754 => 47,            -- (001011.110010 | 11.78125)     => (001.01111 | 1.46875)         
    755 => 47,            -- (001011.110011 | 11.796875)    => (001.01111 | 1.46875)         
    756 => 47,            -- (001011.110100 | 11.8125)      => (001.01111 | 1.46875)         
    757 => 47,            -- (001011.110101 | 11.828125)    => (001.01111 | 1.46875)         
    758 => 47,            -- (001011.110110 | 11.84375)     => (001.01111 | 1.46875)         
    759 => 47,            -- (001011.110111 | 11.859375)    => (001.01111 | 1.46875)         
    760 => 47,            -- (001011.111000 | 11.875)       => (001.01111 | 1.46875)         
    761 => 47,            -- (001011.111001 | 11.890625)    => (001.01111 | 1.46875)         
    762 => 47,            -- (001011.111010 | 11.90625)     => (001.01111 | 1.46875)         
    763 => 47,            -- (001011.111011 | 11.921875)    => (001.01111 | 1.46875)         
    764 => 47,            -- (001011.111100 | 11.9375)      => (001.01111 | 1.46875)         
    765 => 47,            -- (001011.111101 | 11.953125)    => (001.01111 | 1.46875)         
    766 => 47,            -- (001011.111110 | 11.96875)     => (001.01111 | 1.46875)         
    767 => 47,            -- (001011.111111 | 11.984375)    => (001.01111 | 1.46875)         
    768 => 47,            -- (001100.000000 | 12.0)         => (001.01111 | 1.46875)         
    769 => 47,            -- (001100.000001 | 12.015625)    => (001.01111 | 1.46875)         
    770 => 47,            -- (001100.000010 | 12.03125)     => (001.01111 | 1.46875)         
    771 => 47,            -- (001100.000011 | 12.046875)    => (001.01111 | 1.46875)         
    772 => 47,            -- (001100.000100 | 12.0625)      => (001.01111 | 1.46875)         
    773 => 47,            -- (001100.000101 | 12.078125)    => (001.01111 | 1.46875)         
    774 => 47,            -- (001100.000110 | 12.09375)     => (001.01111 | 1.46875)         
    775 => 47,            -- (001100.000111 | 12.109375)    => (001.01111 | 1.46875)         
    776 => 47,            -- (001100.001000 | 12.125)       => (001.01111 | 1.46875)         
    777 => 47,            -- (001100.001001 | 12.140625)    => (001.01111 | 1.46875)         
    778 => 47,            -- (001100.001010 | 12.15625)     => (001.01111 | 1.46875)         
    779 => 47,            -- (001100.001011 | 12.171875)    => (001.01111 | 1.46875)         
    780 => 47,            -- (001100.001100 | 12.1875)      => (001.01111 | 1.46875)         
    781 => 47,            -- (001100.001101 | 12.203125)    => (001.01111 | 1.46875)         
    782 => 47,            -- (001100.001110 | 12.21875)     => (001.01111 | 1.46875)         
    783 => 47,            -- (001100.001111 | 12.234375)    => (001.01111 | 1.46875)         
    784 => 47,            -- (001100.010000 | 12.25)        => (001.01111 | 1.46875)         
    785 => 47,            -- (001100.010001 | 12.265625)    => (001.01111 | 1.46875)         
    786 => 47,            -- (001100.010010 | 12.28125)     => (001.01111 | 1.46875)         
    787 => 47,            -- (001100.010011 | 12.296875)    => (001.01111 | 1.46875)         
    788 => 47,            -- (001100.010100 | 12.3125)      => (001.01111 | 1.46875)         
    789 => 47,            -- (001100.010101 | 12.328125)    => (001.01111 | 1.46875)         
    790 => 47,            -- (001100.010110 | 12.34375)     => (001.01111 | 1.46875)         
    791 => 47,            -- (001100.010111 | 12.359375)    => (001.01111 | 1.46875)         
    792 => 47,            -- (001100.011000 | 12.375)       => (001.01111 | 1.46875)         
    793 => 47,            -- (001100.011001 | 12.390625)    => (001.01111 | 1.46875)         
    794 => 47,            -- (001100.011010 | 12.40625)     => (001.01111 | 1.46875)         
    795 => 47,            -- (001100.011011 | 12.421875)    => (001.01111 | 1.46875)         
    796 => 47,            -- (001100.011100 | 12.4375)      => (001.01111 | 1.46875)         
    797 => 47,            -- (001100.011101 | 12.453125)    => (001.01111 | 1.46875)         
    798 => 47,            -- (001100.011110 | 12.46875)     => (001.01111 | 1.46875)         
    799 => 47,            -- (001100.011111 | 12.484375)    => (001.01111 | 1.46875)         
    800 => 47,            -- (001100.100000 | 12.5)         => (001.01111 | 1.46875)         
    801 => 47,            -- (001100.100001 | 12.515625)    => (001.01111 | 1.46875)         
    802 => 47,            -- (001100.100010 | 12.53125)     => (001.01111 | 1.46875)         
    803 => 47,            -- (001100.100011 | 12.546875)    => (001.01111 | 1.46875)         
    804 => 47,            -- (001100.100100 | 12.5625)      => (001.01111 | 1.46875)         
    805 => 47,            -- (001100.100101 | 12.578125)    => (001.01111 | 1.46875)         
    806 => 47,            -- (001100.100110 | 12.59375)     => (001.01111 | 1.46875)         
    807 => 47,            -- (001100.100111 | 12.609375)    => (001.01111 | 1.46875)         
    808 => 47,            -- (001100.101000 | 12.625)       => (001.01111 | 1.46875)         
    809 => 47,            -- (001100.101001 | 12.640625)    => (001.01111 | 1.46875)         
    810 => 47,            -- (001100.101010 | 12.65625)     => (001.01111 | 1.46875)         
    811 => 47,            -- (001100.101011 | 12.671875)    => (001.01111 | 1.46875)         
    812 => 47,            -- (001100.101100 | 12.6875)      => (001.01111 | 1.46875)         
    813 => 47,            -- (001100.101101 | 12.703125)    => (001.01111 | 1.46875)         
    814 => 47,            -- (001100.101110 | 12.71875)     => (001.01111 | 1.46875)         
    815 => 47,            -- (001100.101111 | 12.734375)    => (001.01111 | 1.46875)         
    816 => 47,            -- (001100.110000 | 12.75)        => (001.01111 | 1.46875)         
    817 => 47,            -- (001100.110001 | 12.765625)    => (001.01111 | 1.46875)         
    818 => 47,            -- (001100.110010 | 12.78125)     => (001.01111 | 1.46875)         
    819 => 47,            -- (001100.110011 | 12.796875)    => (001.01111 | 1.46875)         
    820 => 47,            -- (001100.110100 | 12.8125)      => (001.01111 | 1.46875)         
    821 => 47,            -- (001100.110101 | 12.828125)    => (001.01111 | 1.46875)         
    822 => 47,            -- (001100.110110 | 12.84375)     => (001.01111 | 1.46875)         
    823 => 47,            -- (001100.110111 | 12.859375)    => (001.01111 | 1.46875)         
    824 => 47,            -- (001100.111000 | 12.875)       => (001.01111 | 1.46875)         
    825 => 47,            -- (001100.111001 | 12.890625)    => (001.01111 | 1.46875)         
    826 => 47,            -- (001100.111010 | 12.90625)     => (001.01111 | 1.46875)         
    827 => 47,            -- (001100.111011 | 12.921875)    => (001.01111 | 1.46875)         
    828 => 47,            -- (001100.111100 | 12.9375)      => (001.01111 | 1.46875)         
    829 => 47,            -- (001100.111101 | 12.953125)    => (001.01111 | 1.46875)         
    830 => 47,            -- (001100.111110 | 12.96875)     => (001.01111 | 1.46875)         
    831 => 47,            -- (001100.111111 | 12.984375)    => (001.01111 | 1.46875)         
    832 => 47,            -- (001101.000000 | 13.0)         => (001.01111 | 1.46875)         
    833 => 47,            -- (001101.000001 | 13.015625)    => (001.01111 | 1.46875)         
    834 => 47,            -- (001101.000010 | 13.03125)     => (001.01111 | 1.46875)         
    835 => 47,            -- (001101.000011 | 13.046875)    => (001.01111 | 1.46875)         
    836 => 47,            -- (001101.000100 | 13.0625)      => (001.01111 | 1.46875)         
    837 => 47,            -- (001101.000101 | 13.078125)    => (001.01111 | 1.46875)         
    838 => 47,            -- (001101.000110 | 13.09375)     => (001.01111 | 1.46875)         
    839 => 47,            -- (001101.000111 | 13.109375)    => (001.01111 | 1.46875)         
    840 => 47,            -- (001101.001000 | 13.125)       => (001.01111 | 1.46875)         
    841 => 47,            -- (001101.001001 | 13.140625)    => (001.01111 | 1.46875)         
    842 => 47,            -- (001101.001010 | 13.15625)     => (001.01111 | 1.46875)         
    843 => 47,            -- (001101.001011 | 13.171875)    => (001.01111 | 1.46875)         
    844 => 47,            -- (001101.001100 | 13.1875)      => (001.01111 | 1.46875)         
    845 => 47,            -- (001101.001101 | 13.203125)    => (001.01111 | 1.46875)         
    846 => 47,            -- (001101.001110 | 13.21875)     => (001.01111 | 1.46875)         
    847 => 47,            -- (001101.001111 | 13.234375)    => (001.01111 | 1.46875)         
    848 => 47,            -- (001101.010000 | 13.25)        => (001.01111 | 1.46875)         
    849 => 47,            -- (001101.010001 | 13.265625)    => (001.01111 | 1.46875)         
    850 => 47,            -- (001101.010010 | 13.28125)     => (001.01111 | 1.46875)         
    851 => 47,            -- (001101.010011 | 13.296875)    => (001.01111 | 1.46875)         
    852 => 47,            -- (001101.010100 | 13.3125)      => (001.01111 | 1.46875)         
    853 => 47,            -- (001101.010101 | 13.328125)    => (001.01111 | 1.46875)         
    854 => 47,            -- (001101.010110 | 13.34375)     => (001.01111 | 1.46875)         
    855 => 47,            -- (001101.010111 | 13.359375)    => (001.01111 | 1.46875)         
    856 => 47,            -- (001101.011000 | 13.375)       => (001.01111 | 1.46875)         
    857 => 47,            -- (001101.011001 | 13.390625)    => (001.01111 | 1.46875)         
    858 => 47,            -- (001101.011010 | 13.40625)     => (001.01111 | 1.46875)         
    859 => 47,            -- (001101.011011 | 13.421875)    => (001.01111 | 1.46875)         
    860 => 47,            -- (001101.011100 | 13.4375)      => (001.01111 | 1.46875)         
    861 => 47,            -- (001101.011101 | 13.453125)    => (001.01111 | 1.46875)         
    862 => 47,            -- (001101.011110 | 13.46875)     => (001.01111 | 1.46875)         
    863 => 47,            -- (001101.011111 | 13.484375)    => (001.01111 | 1.46875)         
    864 => 47,            -- (001101.100000 | 13.5)         => (001.01111 | 1.46875)         
    865 => 47,            -- (001101.100001 | 13.515625)    => (001.01111 | 1.46875)         
    866 => 47,            -- (001101.100010 | 13.53125)     => (001.01111 | 1.46875)         
    867 => 47,            -- (001101.100011 | 13.546875)    => (001.01111 | 1.46875)         
    868 => 47,            -- (001101.100100 | 13.5625)      => (001.01111 | 1.46875)         
    869 => 47,            -- (001101.100101 | 13.578125)    => (001.01111 | 1.46875)         
    870 => 47,            -- (001101.100110 | 13.59375)     => (001.01111 | 1.46875)         
    871 => 47,            -- (001101.100111 | 13.609375)    => (001.01111 | 1.46875)         
    872 => 47,            -- (001101.101000 | 13.625)       => (001.01111 | 1.46875)         
    873 => 47,            -- (001101.101001 | 13.640625)    => (001.01111 | 1.46875)         
    874 => 47,            -- (001101.101010 | 13.65625)     => (001.01111 | 1.46875)         
    875 => 47,            -- (001101.101011 | 13.671875)    => (001.01111 | 1.46875)         
    876 => 47,            -- (001101.101100 | 13.6875)      => (001.01111 | 1.46875)         
    877 => 47,            -- (001101.101101 | 13.703125)    => (001.01111 | 1.46875)         
    878 => 47,            -- (001101.101110 | 13.71875)     => (001.01111 | 1.46875)         
    879 => 47,            -- (001101.101111 | 13.734375)    => (001.01111 | 1.46875)         
    880 => 47,            -- (001101.110000 | 13.75)        => (001.01111 | 1.46875)         
    881 => 47,            -- (001101.110001 | 13.765625)    => (001.01111 | 1.46875)         
    882 => 47,            -- (001101.110010 | 13.78125)     => (001.01111 | 1.46875)         
    883 => 47,            -- (001101.110011 | 13.796875)    => (001.01111 | 1.46875)         
    884 => 47,            -- (001101.110100 | 13.8125)      => (001.01111 | 1.46875)         
    885 => 47,            -- (001101.110101 | 13.828125)    => (001.01111 | 1.46875)         
    886 => 47,            -- (001101.110110 | 13.84375)     => (001.01111 | 1.46875)         
    887 => 47,            -- (001101.110111 | 13.859375)    => (001.01111 | 1.46875)         
    888 => 47,            -- (001101.111000 | 13.875)       => (001.01111 | 1.46875)         
    889 => 47,            -- (001101.111001 | 13.890625)    => (001.01111 | 1.46875)         
    890 => 47,            -- (001101.111010 | 13.90625)     => (001.01111 | 1.46875)         
    891 => 47,            -- (001101.111011 | 13.921875)    => (001.01111 | 1.46875)         
    892 => 47,            -- (001101.111100 | 13.9375)      => (001.01111 | 1.46875)         
    893 => 47,            -- (001101.111101 | 13.953125)    => (001.01111 | 1.46875)         
    894 => 47,            -- (001101.111110 | 13.96875)     => (001.01111 | 1.46875)         
    895 => 47,            -- (001101.111111 | 13.984375)    => (001.01111 | 1.46875)         
    896 => 47,            -- (001110.000000 | 14.0)         => (001.01111 | 1.46875)         
    897 => 47,            -- (001110.000001 | 14.015625)    => (001.01111 | 1.46875)         
    898 => 47,            -- (001110.000010 | 14.03125)     => (001.01111 | 1.46875)         
    899 => 47,            -- (001110.000011 | 14.046875)    => (001.01111 | 1.46875)         
    900 => 47,            -- (001110.000100 | 14.0625)      => (001.01111 | 1.46875)         
    901 => 47,            -- (001110.000101 | 14.078125)    => (001.01111 | 1.46875)         
    902 => 47,            -- (001110.000110 | 14.09375)     => (001.01111 | 1.46875)         
    903 => 48,            -- (001110.000111 | 14.109375)    => (001.10000 | 1.5)             
    904 => 48,            -- (001110.001000 | 14.125)       => (001.10000 | 1.5)             
    905 => 48,            -- (001110.001001 | 14.140625)    => (001.10000 | 1.5)             
    906 => 48,            -- (001110.001010 | 14.15625)     => (001.10000 | 1.5)             
    907 => 48,            -- (001110.001011 | 14.171875)    => (001.10000 | 1.5)             
    908 => 48,            -- (001110.001100 | 14.1875)      => (001.10000 | 1.5)             
    909 => 48,            -- (001110.001101 | 14.203125)    => (001.10000 | 1.5)             
    910 => 48,            -- (001110.001110 | 14.21875)     => (001.10000 | 1.5)             
    911 => 48,            -- (001110.001111 | 14.234375)    => (001.10000 | 1.5)             
    912 => 48,            -- (001110.010000 | 14.25)        => (001.10000 | 1.5)             
    913 => 48,            -- (001110.010001 | 14.265625)    => (001.10000 | 1.5)             
    914 => 48,            -- (001110.010010 | 14.28125)     => (001.10000 | 1.5)             
    915 => 48,            -- (001110.010011 | 14.296875)    => (001.10000 | 1.5)             
    916 => 48,            -- (001110.010100 | 14.3125)      => (001.10000 | 1.5)             
    917 => 48,            -- (001110.010101 | 14.328125)    => (001.10000 | 1.5)             
    918 => 48,            -- (001110.010110 | 14.34375)     => (001.10000 | 1.5)             
    919 => 48,            -- (001110.010111 | 14.359375)    => (001.10000 | 1.5)             
    920 => 48,            -- (001110.011000 | 14.375)       => (001.10000 | 1.5)             
    921 => 48,            -- (001110.011001 | 14.390625)    => (001.10000 | 1.5)             
    922 => 48,            -- (001110.011010 | 14.40625)     => (001.10000 | 1.5)             
    923 => 48,            -- (001110.011011 | 14.421875)    => (001.10000 | 1.5)             
    924 => 48,            -- (001110.011100 | 14.4375)      => (001.10000 | 1.5)             
    925 => 48,            -- (001110.011101 | 14.453125)    => (001.10000 | 1.5)             
    926 => 48,            -- (001110.011110 | 14.46875)     => (001.10000 | 1.5)             
    927 => 48,            -- (001110.011111 | 14.484375)    => (001.10000 | 1.5)             
    928 => 48,            -- (001110.100000 | 14.5)         => (001.10000 | 1.5)             
    929 => 48,            -- (001110.100001 | 14.515625)    => (001.10000 | 1.5)             
    930 => 48,            -- (001110.100010 | 14.53125)     => (001.10000 | 1.5)             
    931 => 48,            -- (001110.100011 | 14.546875)    => (001.10000 | 1.5)             
    932 => 48,            -- (001110.100100 | 14.5625)      => (001.10000 | 1.5)             
    933 => 48,            -- (001110.100101 | 14.578125)    => (001.10000 | 1.5)             
    934 => 48,            -- (001110.100110 | 14.59375)     => (001.10000 | 1.5)             
    935 => 48,            -- (001110.100111 | 14.609375)    => (001.10000 | 1.5)             
    936 => 48,            -- (001110.101000 | 14.625)       => (001.10000 | 1.5)             
    937 => 48,            -- (001110.101001 | 14.640625)    => (001.10000 | 1.5)             
    938 => 48,            -- (001110.101010 | 14.65625)     => (001.10000 | 1.5)             
    939 => 48,            -- (001110.101011 | 14.671875)    => (001.10000 | 1.5)             
    940 => 48,            -- (001110.101100 | 14.6875)      => (001.10000 | 1.5)             
    941 => 48,            -- (001110.101101 | 14.703125)    => (001.10000 | 1.5)             
    942 => 48,            -- (001110.101110 | 14.71875)     => (001.10000 | 1.5)             
    943 => 48,            -- (001110.101111 | 14.734375)    => (001.10000 | 1.5)             
    944 => 48,            -- (001110.110000 | 14.75)        => (001.10000 | 1.5)             
    945 => 48,            -- (001110.110001 | 14.765625)    => (001.10000 | 1.5)             
    946 => 48,            -- (001110.110010 | 14.78125)     => (001.10000 | 1.5)             
    947 => 48,            -- (001110.110011 | 14.796875)    => (001.10000 | 1.5)             
    948 => 48,            -- (001110.110100 | 14.8125)      => (001.10000 | 1.5)             
    949 => 48,            -- (001110.110101 | 14.828125)    => (001.10000 | 1.5)             
    950 => 48,            -- (001110.110110 | 14.84375)     => (001.10000 | 1.5)             
    951 => 48,            -- (001110.110111 | 14.859375)    => (001.10000 | 1.5)             
    952 => 48,            -- (001110.111000 | 14.875)       => (001.10000 | 1.5)             
    953 => 48,            -- (001110.111001 | 14.890625)    => (001.10000 | 1.5)             
    954 => 48,            -- (001110.111010 | 14.90625)     => (001.10000 | 1.5)             
    955 => 48,            -- (001110.111011 | 14.921875)    => (001.10000 | 1.5)             
    956 => 48,            -- (001110.111100 | 14.9375)      => (001.10000 | 1.5)             
    957 => 48,            -- (001110.111101 | 14.953125)    => (001.10000 | 1.5)             
    958 => 48,            -- (001110.111110 | 14.96875)     => (001.10000 | 1.5)             
    959 => 48,            -- (001110.111111 | 14.984375)    => (001.10000 | 1.5)             
    960 => 48,            -- (001111.000000 | 15.0)         => (001.10000 | 1.5)             
    961 => 48,            -- (001111.000001 | 15.015625)    => (001.10000 | 1.5)             
    962 => 48,            -- (001111.000010 | 15.03125)     => (001.10000 | 1.5)             
    963 => 48,            -- (001111.000011 | 15.046875)    => (001.10000 | 1.5)             
    964 => 48,            -- (001111.000100 | 15.0625)      => (001.10000 | 1.5)             
    965 => 48,            -- (001111.000101 | 15.078125)    => (001.10000 | 1.5)             
    966 => 48,            -- (001111.000110 | 15.09375)     => (001.10000 | 1.5)             
    967 => 48,            -- (001111.000111 | 15.109375)    => (001.10000 | 1.5)             
    968 => 48,            -- (001111.001000 | 15.125)       => (001.10000 | 1.5)             
    969 => 48,            -- (001111.001001 | 15.140625)    => (001.10000 | 1.5)             
    970 => 48,            -- (001111.001010 | 15.15625)     => (001.10000 | 1.5)             
    971 => 48,            -- (001111.001011 | 15.171875)    => (001.10000 | 1.5)             
    972 => 48,            -- (001111.001100 | 15.1875)      => (001.10000 | 1.5)             
    973 => 48,            -- (001111.001101 | 15.203125)    => (001.10000 | 1.5)             
    974 => 48,            -- (001111.001110 | 15.21875)     => (001.10000 | 1.5)             
    975 => 48,            -- (001111.001111 | 15.234375)    => (001.10000 | 1.5)             
    976 => 48,            -- (001111.010000 | 15.25)        => (001.10000 | 1.5)             
    977 => 48,            -- (001111.010001 | 15.265625)    => (001.10000 | 1.5)             
    978 => 48,            -- (001111.010010 | 15.28125)     => (001.10000 | 1.5)             
    979 => 48,            -- (001111.010011 | 15.296875)    => (001.10000 | 1.5)             
    980 => 48,            -- (001111.010100 | 15.3125)      => (001.10000 | 1.5)             
    981 => 48,            -- (001111.010101 | 15.328125)    => (001.10000 | 1.5)             
    982 => 48,            -- (001111.010110 | 15.34375)     => (001.10000 | 1.5)             
    983 => 48,            -- (001111.010111 | 15.359375)    => (001.10000 | 1.5)             
    984 => 48,            -- (001111.011000 | 15.375)       => (001.10000 | 1.5)             
    985 => 48,            -- (001111.011001 | 15.390625)    => (001.10000 | 1.5)             
    986 => 48,            -- (001111.011010 | 15.40625)     => (001.10000 | 1.5)             
    987 => 48,            -- (001111.011011 | 15.421875)    => (001.10000 | 1.5)             
    988 => 48,            -- (001111.011100 | 15.4375)      => (001.10000 | 1.5)             
    989 => 48,            -- (001111.011101 | 15.453125)    => (001.10000 | 1.5)             
    990 => 48,            -- (001111.011110 | 15.46875)     => (001.10000 | 1.5)             
    991 => 48,            -- (001111.011111 | 15.484375)    => (001.10000 | 1.5)             
    992 => 48,            -- (001111.100000 | 15.5)         => (001.10000 | 1.5)             
    993 => 48,            -- (001111.100001 | 15.515625)    => (001.10000 | 1.5)             
    994 => 48,            -- (001111.100010 | 15.53125)     => (001.10000 | 1.5)             
    995 => 48,            -- (001111.100011 | 15.546875)    => (001.10000 | 1.5)             
    996 => 48,            -- (001111.100100 | 15.5625)      => (001.10000 | 1.5)             
    997 => 48,            -- (001111.100101 | 15.578125)    => (001.10000 | 1.5)             
    998 => 48,            -- (001111.100110 | 15.59375)     => (001.10000 | 1.5)             
    999 => 48,            -- (001111.100111 | 15.609375)    => (001.10000 | 1.5)             
    1000 => 48,           -- (001111.101000 | 15.625)       => (001.10000 | 1.5)             
    1001 => 48,           -- (001111.101001 | 15.640625)    => (001.10000 | 1.5)             
    1002 => 48,           -- (001111.101010 | 15.65625)     => (001.10000 | 1.5)             
    1003 => 48,           -- (001111.101011 | 15.671875)    => (001.10000 | 1.5)             
    1004 => 48,           -- (001111.101100 | 15.6875)      => (001.10000 | 1.5)             
    1005 => 48,           -- (001111.101101 | 15.703125)    => (001.10000 | 1.5)             
    1006 => 48,           -- (001111.101110 | 15.71875)     => (001.10000 | 1.5)             
    1007 => 48,           -- (001111.101111 | 15.734375)    => (001.10000 | 1.5)             
    1008 => 48,           -- (001111.110000 | 15.75)        => (001.10000 | 1.5)             
    1009 => 48,           -- (001111.110001 | 15.765625)    => (001.10000 | 1.5)             
    1010 => 48,           -- (001111.110010 | 15.78125)     => (001.10000 | 1.5)             
    1011 => 48,           -- (001111.110011 | 15.796875)    => (001.10000 | 1.5)             
    1012 => 48,           -- (001111.110100 | 15.8125)      => (001.10000 | 1.5)             
    1013 => 48,           -- (001111.110101 | 15.828125)    => (001.10000 | 1.5)             
    1014 => 48,           -- (001111.110110 | 15.84375)     => (001.10000 | 1.5)             
    1015 => 48,           -- (001111.110111 | 15.859375)    => (001.10000 | 1.5)             
    1016 => 48,           -- (001111.111000 | 15.875)       => (001.10000 | 1.5)             
    1017 => 48,           -- (001111.111001 | 15.890625)    => (001.10000 | 1.5)             
    1018 => 48,           -- (001111.111010 | 15.90625)     => (001.10000 | 1.5)             
    1019 => 48,           -- (001111.111011 | 15.921875)    => (001.10000 | 1.5)             
    1020 => 48,           -- (001111.111100 | 15.9375)      => (001.10000 | 1.5)             
    1021 => 48,           -- (001111.111101 | 15.953125)    => (001.10000 | 1.5)             
    1022 => 48,           -- (001111.111110 | 15.96875)     => (001.10000 | 1.5)             
    1023 => 48,           -- (001111.111111 | 15.984375)    => (001.10000 | 1.5)             
    1024 => 48,           -- (010000.000000 | 16.0)         => (001.10000 | 1.5)             
    1025 => 48,           -- (010000.000001 | 16.015625)    => (001.10000 | 1.5)             
    1026 => 48,           -- (010000.000010 | 16.03125)     => (001.10000 | 1.5)             
    1027 => 48,           -- (010000.000011 | 16.046875)    => (001.10000 | 1.5)             
    1028 => 48,           -- (010000.000100 | 16.0625)      => (001.10000 | 1.5)             
    1029 => 48,           -- (010000.000101 | 16.078125)    => (001.10000 | 1.5)             
    1030 => 48,           -- (010000.000110 | 16.09375)     => (001.10000 | 1.5)             
    1031 => 48,           -- (010000.000111 | 16.109375)    => (001.10000 | 1.5)             
    1032 => 48,           -- (010000.001000 | 16.125)       => (001.10000 | 1.5)             
    1033 => 48,           -- (010000.001001 | 16.140625)    => (001.10000 | 1.5)             
    1034 => 48,           -- (010000.001010 | 16.15625)     => (001.10000 | 1.5)             
    1035 => 48,           -- (010000.001011 | 16.171875)    => (001.10000 | 1.5)             
    1036 => 48,           -- (010000.001100 | 16.1875)      => (001.10000 | 1.5)             
    1037 => 48,           -- (010000.001101 | 16.203125)    => (001.10000 | 1.5)             
    1038 => 48,           -- (010000.001110 | 16.21875)     => (001.10000 | 1.5)             
    1039 => 48,           -- (010000.001111 | 16.234375)    => (001.10000 | 1.5)             
    1040 => 48,           -- (010000.010000 | 16.25)        => (001.10000 | 1.5)             
    1041 => 48,           -- (010000.010001 | 16.265625)    => (001.10000 | 1.5)             
    1042 => 48,           -- (010000.010010 | 16.28125)     => (001.10000 | 1.5)             
    1043 => 48,           -- (010000.010011 | 16.296875)    => (001.10000 | 1.5)             
    1044 => 48,           -- (010000.010100 | 16.3125)      => (001.10000 | 1.5)             
    1045 => 48,           -- (010000.010101 | 16.328125)    => (001.10000 | 1.5)             
    1046 => 48,           -- (010000.010110 | 16.34375)     => (001.10000 | 1.5)             
    1047 => 48,           -- (010000.010111 | 16.359375)    => (001.10000 | 1.5)             
    1048 => 48,           -- (010000.011000 | 16.375)       => (001.10000 | 1.5)             
    1049 => 48,           -- (010000.011001 | 16.390625)    => (001.10000 | 1.5)             
    1050 => 48,           -- (010000.011010 | 16.40625)     => (001.10000 | 1.5)             
    1051 => 48,           -- (010000.011011 | 16.421875)    => (001.10000 | 1.5)             
    1052 => 48,           -- (010000.011100 | 16.4375)      => (001.10000 | 1.5)             
    1053 => 48,           -- (010000.011101 | 16.453125)    => (001.10000 | 1.5)             
    1054 => 48,           -- (010000.011110 | 16.46875)     => (001.10000 | 1.5)             
    1055 => 48,           -- (010000.011111 | 16.484375)    => (001.10000 | 1.5)             
    1056 => 48,           -- (010000.100000 | 16.5)         => (001.10000 | 1.5)             
    1057 => 48,           -- (010000.100001 | 16.515625)    => (001.10000 | 1.5)             
    1058 => 48,           -- (010000.100010 | 16.53125)     => (001.10000 | 1.5)             
    1059 => 48,           -- (010000.100011 | 16.546875)    => (001.10000 | 1.5)             
    1060 => 48,           -- (010000.100100 | 16.5625)      => (001.10000 | 1.5)             
    1061 => 48,           -- (010000.100101 | 16.578125)    => (001.10000 | 1.5)             
    1062 => 48,           -- (010000.100110 | 16.59375)     => (001.10000 | 1.5)             
    1063 => 48,           -- (010000.100111 | 16.609375)    => (001.10000 | 1.5)             
    1064 => 48,           -- (010000.101000 | 16.625)       => (001.10000 | 1.5)             
    1065 => 48,           -- (010000.101001 | 16.640625)    => (001.10000 | 1.5)             
    1066 => 48,           -- (010000.101010 | 16.65625)     => (001.10000 | 1.5)             
    1067 => 48,           -- (010000.101011 | 16.671875)    => (001.10000 | 1.5)             
    1068 => 48,           -- (010000.101100 | 16.6875)      => (001.10000 | 1.5)             
    1069 => 48,           -- (010000.101101 | 16.703125)    => (001.10000 | 1.5)             
    1070 => 48,           -- (010000.101110 | 16.71875)     => (001.10000 | 1.5)             
    1071 => 48,           -- (010000.101111 | 16.734375)    => (001.10000 | 1.5)             
    1072 => 48,           -- (010000.110000 | 16.75)        => (001.10000 | 1.5)             
    1073 => 48,           -- (010000.110001 | 16.765625)    => (001.10000 | 1.5)             
    1074 => 48,           -- (010000.110010 | 16.78125)     => (001.10000 | 1.5)             
    1075 => 48,           -- (010000.110011 | 16.796875)    => (001.10000 | 1.5)             
    1076 => 48,           -- (010000.110100 | 16.8125)      => (001.10000 | 1.5)             
    1077 => 48,           -- (010000.110101 | 16.828125)    => (001.10000 | 1.5)             
    1078 => 48,           -- (010000.110110 | 16.84375)     => (001.10000 | 1.5)             
    1079 => 48,           -- (010000.110111 | 16.859375)    => (001.10000 | 1.5)             
    1080 => 48,           -- (010000.111000 | 16.875)       => (001.10000 | 1.5)             
    1081 => 48,           -- (010000.111001 | 16.890625)    => (001.10000 | 1.5)             
    1082 => 48,           -- (010000.111010 | 16.90625)     => (001.10000 | 1.5)             
    1083 => 48,           -- (010000.111011 | 16.921875)    => (001.10000 | 1.5)             
    1084 => 48,           -- (010000.111100 | 16.9375)      => (001.10000 | 1.5)             
    1085 => 48,           -- (010000.111101 | 16.953125)    => (001.10000 | 1.5)             
    1086 => 48,           -- (010000.111110 | 16.96875)     => (001.10000 | 1.5)             
    1087 => 48,           -- (010000.111111 | 16.984375)    => (001.10000 | 1.5)             
    1088 => 48,           -- (010001.000000 | 17.0)         => (001.10000 | 1.5)             
    1089 => 48,           -- (010001.000001 | 17.015625)    => (001.10000 | 1.5)             
    1090 => 48,           -- (010001.000010 | 17.03125)     => (001.10000 | 1.5)             
    1091 => 48,           -- (010001.000011 | 17.046875)    => (001.10000 | 1.5)             
    1092 => 48,           -- (010001.000100 | 17.0625)      => (001.10000 | 1.5)             
    1093 => 48,           -- (010001.000101 | 17.078125)    => (001.10000 | 1.5)             
    1094 => 48,           -- (010001.000110 | 17.09375)     => (001.10000 | 1.5)             
    1095 => 48,           -- (010001.000111 | 17.109375)    => (001.10000 | 1.5)             
    1096 => 48,           -- (010001.001000 | 17.125)       => (001.10000 | 1.5)             
    1097 => 48,           -- (010001.001001 | 17.140625)    => (001.10000 | 1.5)             
    1098 => 48,           -- (010001.001010 | 17.15625)     => (001.10000 | 1.5)             
    1099 => 48,           -- (010001.001011 | 17.171875)    => (001.10000 | 1.5)             
    1100 => 48,           -- (010001.001100 | 17.1875)      => (001.10000 | 1.5)             
    1101 => 48,           -- (010001.001101 | 17.203125)    => (001.10000 | 1.5)             
    1102 => 48,           -- (010001.001110 | 17.21875)     => (001.10000 | 1.5)             
    1103 => 48,           -- (010001.001111 | 17.234375)    => (001.10000 | 1.5)             
    1104 => 48,           -- (010001.010000 | 17.25)        => (001.10000 | 1.5)             
    1105 => 48,           -- (010001.010001 | 17.265625)    => (001.10000 | 1.5)             
    1106 => 48,           -- (010001.010010 | 17.28125)     => (001.10000 | 1.5)             
    1107 => 48,           -- (010001.010011 | 17.296875)    => (001.10000 | 1.5)             
    1108 => 48,           -- (010001.010100 | 17.3125)      => (001.10000 | 1.5)             
    1109 => 48,           -- (010001.010101 | 17.328125)    => (001.10000 | 1.5)             
    1110 => 48,           -- (010001.010110 | 17.34375)     => (001.10000 | 1.5)             
    1111 => 48,           -- (010001.010111 | 17.359375)    => (001.10000 | 1.5)             
    1112 => 48,           -- (010001.011000 | 17.375)       => (001.10000 | 1.5)             
    1113 => 48,           -- (010001.011001 | 17.390625)    => (001.10000 | 1.5)             
    1114 => 48,           -- (010001.011010 | 17.40625)     => (001.10000 | 1.5)             
    1115 => 48,           -- (010001.011011 | 17.421875)    => (001.10000 | 1.5)             
    1116 => 48,           -- (010001.011100 | 17.4375)      => (001.10000 | 1.5)             
    1117 => 48,           -- (010001.011101 | 17.453125)    => (001.10000 | 1.5)             
    1118 => 48,           -- (010001.011110 | 17.46875)     => (001.10000 | 1.5)             
    1119 => 48,           -- (010001.011111 | 17.484375)    => (001.10000 | 1.5)             
    1120 => 48,           -- (010001.100000 | 17.5)         => (001.10000 | 1.5)             
    1121 => 48,           -- (010001.100001 | 17.515625)    => (001.10000 | 1.5)             
    1122 => 48,           -- (010001.100010 | 17.53125)     => (001.10000 | 1.5)             
    1123 => 48,           -- (010001.100011 | 17.546875)    => (001.10000 | 1.5)             
    1124 => 48,           -- (010001.100100 | 17.5625)      => (001.10000 | 1.5)             
    1125 => 48,           -- (010001.100101 | 17.578125)    => (001.10000 | 1.5)             
    1126 => 48,           -- (010001.100110 | 17.59375)     => (001.10000 | 1.5)             
    1127 => 48,           -- (010001.100111 | 17.609375)    => (001.10000 | 1.5)             
    1128 => 48,           -- (010001.101000 | 17.625)       => (001.10000 | 1.5)             
    1129 => 48,           -- (010001.101001 | 17.640625)    => (001.10000 | 1.5)             
    1130 => 48,           -- (010001.101010 | 17.65625)     => (001.10000 | 1.5)             
    1131 => 48,           -- (010001.101011 | 17.671875)    => (001.10000 | 1.5)             
    1132 => 48,           -- (010001.101100 | 17.6875)      => (001.10000 | 1.5)             
    1133 => 48,           -- (010001.101101 | 17.703125)    => (001.10000 | 1.5)             
    1134 => 48,           -- (010001.101110 | 17.71875)     => (001.10000 | 1.5)             
    1135 => 48,           -- (010001.101111 | 17.734375)    => (001.10000 | 1.5)             
    1136 => 48,           -- (010001.110000 | 17.75)        => (001.10000 | 1.5)             
    1137 => 48,           -- (010001.110001 | 17.765625)    => (001.10000 | 1.5)             
    1138 => 48,           -- (010001.110010 | 17.78125)     => (001.10000 | 1.5)             
    1139 => 48,           -- (010001.110011 | 17.796875)    => (001.10000 | 1.5)             
    1140 => 48,           -- (010001.110100 | 17.8125)      => (001.10000 | 1.5)             
    1141 => 48,           -- (010001.110101 | 17.828125)    => (001.10000 | 1.5)             
    1142 => 48,           -- (010001.110110 | 17.84375)     => (001.10000 | 1.5)             
    1143 => 48,           -- (010001.110111 | 17.859375)    => (001.10000 | 1.5)             
    1144 => 48,           -- (010001.111000 | 17.875)       => (001.10000 | 1.5)             
    1145 => 48,           -- (010001.111001 | 17.890625)    => (001.10000 | 1.5)             
    1146 => 48,           -- (010001.111010 | 17.90625)     => (001.10000 | 1.5)             
    1147 => 48,           -- (010001.111011 | 17.921875)    => (001.10000 | 1.5)             
    1148 => 48,           -- (010001.111100 | 17.9375)      => (001.10000 | 1.5)             
    1149 => 48,           -- (010001.111101 | 17.953125)    => (001.10000 | 1.5)             
    1150 => 48,           -- (010001.111110 | 17.96875)     => (001.10000 | 1.5)             
    1151 => 48,           -- (010001.111111 | 17.984375)    => (001.10000 | 1.5)             
    1152 => 48,           -- (010010.000000 | 18.0)         => (001.10000 | 1.5)             
    1153 => 48,           -- (010010.000001 | 18.015625)    => (001.10000 | 1.5)             
    1154 => 48,           -- (010010.000010 | 18.03125)     => (001.10000 | 1.5)             
    1155 => 48,           -- (010010.000011 | 18.046875)    => (001.10000 | 1.5)             
    1156 => 48,           -- (010010.000100 | 18.0625)      => (001.10000 | 1.5)             
    1157 => 48,           -- (010010.000101 | 18.078125)    => (001.10000 | 1.5)             
    1158 => 48,           -- (010010.000110 | 18.09375)     => (001.10000 | 1.5)             
    1159 => 48,           -- (010010.000111 | 18.109375)    => (001.10000 | 1.5)             
    1160 => 48,           -- (010010.001000 | 18.125)       => (001.10000 | 1.5)             
    1161 => 48,           -- (010010.001001 | 18.140625)    => (001.10000 | 1.5)             
    1162 => 48,           -- (010010.001010 | 18.15625)     => (001.10000 | 1.5)             
    1163 => 48,           -- (010010.001011 | 18.171875)    => (001.10000 | 1.5)             
    1164 => 48,           -- (010010.001100 | 18.1875)      => (001.10000 | 1.5)             
    1165 => 48,           -- (010010.001101 | 18.203125)    => (001.10000 | 1.5)             
    1166 => 48,           -- (010010.001110 | 18.21875)     => (001.10000 | 1.5)             
    1167 => 48,           -- (010010.001111 | 18.234375)    => (001.10000 | 1.5)             
    1168 => 48,           -- (010010.010000 | 18.25)        => (001.10000 | 1.5)             
    1169 => 48,           -- (010010.010001 | 18.265625)    => (001.10000 | 1.5)             
    1170 => 48,           -- (010010.010010 | 18.28125)     => (001.10000 | 1.5)             
    1171 => 48,           -- (010010.010011 | 18.296875)    => (001.10000 | 1.5)             
    1172 => 48,           -- (010010.010100 | 18.3125)      => (001.10000 | 1.5)             
    1173 => 48,           -- (010010.010101 | 18.328125)    => (001.10000 | 1.5)             
    1174 => 48,           -- (010010.010110 | 18.34375)     => (001.10000 | 1.5)             
    1175 => 48,           -- (010010.010111 | 18.359375)    => (001.10000 | 1.5)             
    1176 => 48,           -- (010010.011000 | 18.375)       => (001.10000 | 1.5)             
    1177 => 48,           -- (010010.011001 | 18.390625)    => (001.10000 | 1.5)             
    1178 => 48,           -- (010010.011010 | 18.40625)     => (001.10000 | 1.5)             
    1179 => 48,           -- (010010.011011 | 18.421875)    => (001.10000 | 1.5)             
    1180 => 48,           -- (010010.011100 | 18.4375)      => (001.10000 | 1.5)             
    1181 => 48,           -- (010010.011101 | 18.453125)    => (001.10000 | 1.5)             
    1182 => 48,           -- (010010.011110 | 18.46875)     => (001.10000 | 1.5)             
    1183 => 48,           -- (010010.011111 | 18.484375)    => (001.10000 | 1.5)             
    1184 => 48,           -- (010010.100000 | 18.5)         => (001.10000 | 1.5)             
    1185 => 48,           -- (010010.100001 | 18.515625)    => (001.10000 | 1.5)             
    1186 => 48,           -- (010010.100010 | 18.53125)     => (001.10000 | 1.5)             
    1187 => 48,           -- (010010.100011 | 18.546875)    => (001.10000 | 1.5)             
    1188 => 48,           -- (010010.100100 | 18.5625)      => (001.10000 | 1.5)             
    1189 => 48,           -- (010010.100101 | 18.578125)    => (001.10000 | 1.5)             
    1190 => 48,           -- (010010.100110 | 18.59375)     => (001.10000 | 1.5)             
    1191 => 48,           -- (010010.100111 | 18.609375)    => (001.10000 | 1.5)             
    1192 => 48,           -- (010010.101000 | 18.625)       => (001.10000 | 1.5)             
    1193 => 48,           -- (010010.101001 | 18.640625)    => (001.10000 | 1.5)             
    1194 => 48,           -- (010010.101010 | 18.65625)     => (001.10000 | 1.5)             
    1195 => 48,           -- (010010.101011 | 18.671875)    => (001.10000 | 1.5)             
    1196 => 48,           -- (010010.101100 | 18.6875)      => (001.10000 | 1.5)             
    1197 => 48,           -- (010010.101101 | 18.703125)    => (001.10000 | 1.5)             
    1198 => 48,           -- (010010.101110 | 18.71875)     => (001.10000 | 1.5)             
    1199 => 48,           -- (010010.101111 | 18.734375)    => (001.10000 | 1.5)             
    1200 => 48,           -- (010010.110000 | 18.75)        => (001.10000 | 1.5)             
    1201 => 48,           -- (010010.110001 | 18.765625)    => (001.10000 | 1.5)             
    1202 => 48,           -- (010010.110010 | 18.78125)     => (001.10000 | 1.5)             
    1203 => 48,           -- (010010.110011 | 18.796875)    => (001.10000 | 1.5)             
    1204 => 48,           -- (010010.110100 | 18.8125)      => (001.10000 | 1.5)             
    1205 => 48,           -- (010010.110101 | 18.828125)    => (001.10000 | 1.5)             
    1206 => 48,           -- (010010.110110 | 18.84375)     => (001.10000 | 1.5)             
    1207 => 48,           -- (010010.110111 | 18.859375)    => (001.10000 | 1.5)             
    1208 => 48,           -- (010010.111000 | 18.875)       => (001.10000 | 1.5)             
    1209 => 48,           -- (010010.111001 | 18.890625)    => (001.10000 | 1.5)             
    1210 => 48,           -- (010010.111010 | 18.90625)     => (001.10000 | 1.5)             
    1211 => 48,           -- (010010.111011 | 18.921875)    => (001.10000 | 1.5)             
    1212 => 48,           -- (010010.111100 | 18.9375)      => (001.10000 | 1.5)             
    1213 => 48,           -- (010010.111101 | 18.953125)    => (001.10000 | 1.5)             
    1214 => 48,           -- (010010.111110 | 18.96875)     => (001.10000 | 1.5)             
    1215 => 48,           -- (010010.111111 | 18.984375)    => (001.10000 | 1.5)             
    1216 => 48,           -- (010011.000000 | 19.0)         => (001.10000 | 1.5)             
    1217 => 48,           -- (010011.000001 | 19.015625)    => (001.10000 | 1.5)             
    1218 => 48,           -- (010011.000010 | 19.03125)     => (001.10000 | 1.5)             
    1219 => 48,           -- (010011.000011 | 19.046875)    => (001.10000 | 1.5)             
    1220 => 48,           -- (010011.000100 | 19.0625)      => (001.10000 | 1.5)             
    1221 => 48,           -- (010011.000101 | 19.078125)    => (001.10000 | 1.5)             
    1222 => 48,           -- (010011.000110 | 19.09375)     => (001.10000 | 1.5)             
    1223 => 48,           -- (010011.000111 | 19.109375)    => (001.10000 | 1.5)             
    1224 => 48,           -- (010011.001000 | 19.125)       => (001.10000 | 1.5)             
    1225 => 48,           -- (010011.001001 | 19.140625)    => (001.10000 | 1.5)             
    1226 => 48,           -- (010011.001010 | 19.15625)     => (001.10000 | 1.5)             
    1227 => 48,           -- (010011.001011 | 19.171875)    => (001.10000 | 1.5)             
    1228 => 48,           -- (010011.001100 | 19.1875)      => (001.10000 | 1.5)             
    1229 => 48,           -- (010011.001101 | 19.203125)    => (001.10000 | 1.5)             
    1230 => 48,           -- (010011.001110 | 19.21875)     => (001.10000 | 1.5)             
    1231 => 48,           -- (010011.001111 | 19.234375)    => (001.10000 | 1.5)             
    1232 => 48,           -- (010011.010000 | 19.25)        => (001.10000 | 1.5)             
    1233 => 48,           -- (010011.010001 | 19.265625)    => (001.10000 | 1.5)             
    1234 => 48,           -- (010011.010010 | 19.28125)     => (001.10000 | 1.5)             
    1235 => 48,           -- (010011.010011 | 19.296875)    => (001.10000 | 1.5)             
    1236 => 48,           -- (010011.010100 | 19.3125)      => (001.10000 | 1.5)             
    1237 => 48,           -- (010011.010101 | 19.328125)    => (001.10000 | 1.5)             
    1238 => 48,           -- (010011.010110 | 19.34375)     => (001.10000 | 1.5)             
    1239 => 48,           -- (010011.010111 | 19.359375)    => (001.10000 | 1.5)             
    1240 => 48,           -- (010011.011000 | 19.375)       => (001.10000 | 1.5)             
    1241 => 48,           -- (010011.011001 | 19.390625)    => (001.10000 | 1.5)             
    1242 => 48,           -- (010011.011010 | 19.40625)     => (001.10000 | 1.5)             
    1243 => 48,           -- (010011.011011 | 19.421875)    => (001.10000 | 1.5)             
    1244 => 48,           -- (010011.011100 | 19.4375)      => (001.10000 | 1.5)             
    1245 => 48,           -- (010011.011101 | 19.453125)    => (001.10000 | 1.5)             
    1246 => 48,           -- (010011.011110 | 19.46875)     => (001.10000 | 1.5)             
    1247 => 48,           -- (010011.011111 | 19.484375)    => (001.10000 | 1.5)             
    1248 => 48,           -- (010011.100000 | 19.5)         => (001.10000 | 1.5)             
    1249 => 48,           -- (010011.100001 | 19.515625)    => (001.10000 | 1.5)             
    1250 => 48,           -- (010011.100010 | 19.53125)     => (001.10000 | 1.5)             
    1251 => 48,           -- (010011.100011 | 19.546875)    => (001.10000 | 1.5)             
    1252 => 48,           -- (010011.100100 | 19.5625)      => (001.10000 | 1.5)             
    1253 => 48,           -- (010011.100101 | 19.578125)    => (001.10000 | 1.5)             
    1254 => 48,           -- (010011.100110 | 19.59375)     => (001.10000 | 1.5)             
    1255 => 48,           -- (010011.100111 | 19.609375)    => (001.10000 | 1.5)             
    1256 => 48,           -- (010011.101000 | 19.625)       => (001.10000 | 1.5)             
    1257 => 48,           -- (010011.101001 | 19.640625)    => (001.10000 | 1.5)             
    1258 => 48,           -- (010011.101010 | 19.65625)     => (001.10000 | 1.5)             
    1259 => 48,           -- (010011.101011 | 19.671875)    => (001.10000 | 1.5)             
    1260 => 48,           -- (010011.101100 | 19.6875)      => (001.10000 | 1.5)             
    1261 => 48,           -- (010011.101101 | 19.703125)    => (001.10000 | 1.5)             
    1262 => 48,           -- (010011.101110 | 19.71875)     => (001.10000 | 1.5)             
    1263 => 48,           -- (010011.101111 | 19.734375)    => (001.10000 | 1.5)             
    1264 => 48,           -- (010011.110000 | 19.75)        => (001.10000 | 1.5)             
    1265 => 48,           -- (010011.110001 | 19.765625)    => (001.10000 | 1.5)             
    1266 => 48,           -- (010011.110010 | 19.78125)     => (001.10000 | 1.5)             
    1267 => 48,           -- (010011.110011 | 19.796875)    => (001.10000 | 1.5)             
    1268 => 48,           -- (010011.110100 | 19.8125)      => (001.10000 | 1.5)             
    1269 => 48,           -- (010011.110101 | 19.828125)    => (001.10000 | 1.5)             
    1270 => 48,           -- (010011.110110 | 19.84375)     => (001.10000 | 1.5)             
    1271 => 48,           -- (010011.110111 | 19.859375)    => (001.10000 | 1.5)             
    1272 => 48,           -- (010011.111000 | 19.875)       => (001.10000 | 1.5)             
    1273 => 48,           -- (010011.111001 | 19.890625)    => (001.10000 | 1.5)             
    1274 => 48,           -- (010011.111010 | 19.90625)     => (001.10000 | 1.5)             
    1275 => 48,           -- (010011.111011 | 19.921875)    => (001.10000 | 1.5)             
    1276 => 48,           -- (010011.111100 | 19.9375)      => (001.10000 | 1.5)             
    1277 => 48,           -- (010011.111101 | 19.953125)    => (001.10000 | 1.5)             
    1278 => 48,           -- (010011.111110 | 19.96875)     => (001.10000 | 1.5)             
    1279 => 48,           -- (010011.111111 | 19.984375)    => (001.10000 | 1.5)             
    1280 => 48,           -- (010100.000000 | 20.0)         => (001.10000 | 1.5)             
    1281 => 48,           -- (010100.000001 | 20.015625)    => (001.10000 | 1.5)             
    1282 => 48,           -- (010100.000010 | 20.03125)     => (001.10000 | 1.5)             
    1283 => 48,           -- (010100.000011 | 20.046875)    => (001.10000 | 1.5)             
    1284 => 48,           -- (010100.000100 | 20.0625)      => (001.10000 | 1.5)             
    1285 => 48,           -- (010100.000101 | 20.078125)    => (001.10000 | 1.5)             
    1286 => 48,           -- (010100.000110 | 20.09375)     => (001.10000 | 1.5)             
    1287 => 48,           -- (010100.000111 | 20.109375)    => (001.10000 | 1.5)             
    1288 => 48,           -- (010100.001000 | 20.125)       => (001.10000 | 1.5)             
    1289 => 48,           -- (010100.001001 | 20.140625)    => (001.10000 | 1.5)             
    1290 => 48,           -- (010100.001010 | 20.15625)     => (001.10000 | 1.5)             
    1291 => 48,           -- (010100.001011 | 20.171875)    => (001.10000 | 1.5)             
    1292 => 48,           -- (010100.001100 | 20.1875)      => (001.10000 | 1.5)             
    1293 => 48,           -- (010100.001101 | 20.203125)    => (001.10000 | 1.5)             
    1294 => 48,           -- (010100.001110 | 20.21875)     => (001.10000 | 1.5)             
    1295 => 48,           -- (010100.001111 | 20.234375)    => (001.10000 | 1.5)             
    1296 => 48,           -- (010100.010000 | 20.25)        => (001.10000 | 1.5)             
    1297 => 48,           -- (010100.010001 | 20.265625)    => (001.10000 | 1.5)             
    1298 => 48,           -- (010100.010010 | 20.28125)     => (001.10000 | 1.5)             
    1299 => 48,           -- (010100.010011 | 20.296875)    => (001.10000 | 1.5)             
    1300 => 48,           -- (010100.010100 | 20.3125)      => (001.10000 | 1.5)             
    1301 => 48,           -- (010100.010101 | 20.328125)    => (001.10000 | 1.5)             
    1302 => 48,           -- (010100.010110 | 20.34375)     => (001.10000 | 1.5)             
    1303 => 48,           -- (010100.010111 | 20.359375)    => (001.10000 | 1.5)             
    1304 => 48,           -- (010100.011000 | 20.375)       => (001.10000 | 1.5)             
    1305 => 48,           -- (010100.011001 | 20.390625)    => (001.10000 | 1.5)             
    1306 => 48,           -- (010100.011010 | 20.40625)     => (001.10000 | 1.5)             
    1307 => 48,           -- (010100.011011 | 20.421875)    => (001.10000 | 1.5)             
    1308 => 48,           -- (010100.011100 | 20.4375)      => (001.10000 | 1.5)             
    1309 => 48,           -- (010100.011101 | 20.453125)    => (001.10000 | 1.5)             
    1310 => 48,           -- (010100.011110 | 20.46875)     => (001.10000 | 1.5)             
    1311 => 48,           -- (010100.011111 | 20.484375)    => (001.10000 | 1.5)             
    1312 => 48,           -- (010100.100000 | 20.5)         => (001.10000 | 1.5)             
    1313 => 48,           -- (010100.100001 | 20.515625)    => (001.10000 | 1.5)             
    1314 => 48,           -- (010100.100010 | 20.53125)     => (001.10000 | 1.5)             
    1315 => 48,           -- (010100.100011 | 20.546875)    => (001.10000 | 1.5)             
    1316 => 48,           -- (010100.100100 | 20.5625)      => (001.10000 | 1.5)             
    1317 => 48,           -- (010100.100101 | 20.578125)    => (001.10000 | 1.5)             
    1318 => 48,           -- (010100.100110 | 20.59375)     => (001.10000 | 1.5)             
    1319 => 48,           -- (010100.100111 | 20.609375)    => (001.10000 | 1.5)             
    1320 => 48,           -- (010100.101000 | 20.625)       => (001.10000 | 1.5)             
    1321 => 48,           -- (010100.101001 | 20.640625)    => (001.10000 | 1.5)             
    1322 => 48,           -- (010100.101010 | 20.65625)     => (001.10000 | 1.5)             
    1323 => 48,           -- (010100.101011 | 20.671875)    => (001.10000 | 1.5)             
    1324 => 48,           -- (010100.101100 | 20.6875)      => (001.10000 | 1.5)             
    1325 => 48,           -- (010100.101101 | 20.703125)    => (001.10000 | 1.5)             
    1326 => 48,           -- (010100.101110 | 20.71875)     => (001.10000 | 1.5)             
    1327 => 48,           -- (010100.101111 | 20.734375)    => (001.10000 | 1.5)             
    1328 => 48,           -- (010100.110000 | 20.75)        => (001.10000 | 1.5)             
    1329 => 48,           -- (010100.110001 | 20.765625)    => (001.10000 | 1.5)             
    1330 => 48,           -- (010100.110010 | 20.78125)     => (001.10000 | 1.5)             
    1331 => 48,           -- (010100.110011 | 20.796875)    => (001.10000 | 1.5)             
    1332 => 48,           -- (010100.110100 | 20.8125)      => (001.10000 | 1.5)             
    1333 => 48,           -- (010100.110101 | 20.828125)    => (001.10000 | 1.5)             
    1334 => 48,           -- (010100.110110 | 20.84375)     => (001.10000 | 1.5)             
    1335 => 48,           -- (010100.110111 | 20.859375)    => (001.10000 | 1.5)             
    1336 => 48,           -- (010100.111000 | 20.875)       => (001.10000 | 1.5)             
    1337 => 48,           -- (010100.111001 | 20.890625)    => (001.10000 | 1.5)             
    1338 => 48,           -- (010100.111010 | 20.90625)     => (001.10000 | 1.5)             
    1339 => 48,           -- (010100.111011 | 20.921875)    => (001.10000 | 1.5)             
    1340 => 48,           -- (010100.111100 | 20.9375)      => (001.10000 | 1.5)             
    1341 => 48,           -- (010100.111101 | 20.953125)    => (001.10000 | 1.5)             
    1342 => 48,           -- (010100.111110 | 20.96875)     => (001.10000 | 1.5)             
    1343 => 48,           -- (010100.111111 | 20.984375)    => (001.10000 | 1.5)             
    1344 => 48,           -- (010101.000000 | 21.0)         => (001.10000 | 1.5)             
    1345 => 48,           -- (010101.000001 | 21.015625)    => (001.10000 | 1.5)             
    1346 => 48,           -- (010101.000010 | 21.03125)     => (001.10000 | 1.5)             
    1347 => 48,           -- (010101.000011 | 21.046875)    => (001.10000 | 1.5)             
    1348 => 48,           -- (010101.000100 | 21.0625)      => (001.10000 | 1.5)             
    1349 => 48,           -- (010101.000101 | 21.078125)    => (001.10000 | 1.5)             
    1350 => 48,           -- (010101.000110 | 21.09375)     => (001.10000 | 1.5)             
    1351 => 48,           -- (010101.000111 | 21.109375)    => (001.10000 | 1.5)             
    1352 => 48,           -- (010101.001000 | 21.125)       => (001.10000 | 1.5)             
    1353 => 48,           -- (010101.001001 | 21.140625)    => (001.10000 | 1.5)             
    1354 => 48,           -- (010101.001010 | 21.15625)     => (001.10000 | 1.5)             
    1355 => 48,           -- (010101.001011 | 21.171875)    => (001.10000 | 1.5)             
    1356 => 48,           -- (010101.001100 | 21.1875)      => (001.10000 | 1.5)             
    1357 => 48,           -- (010101.001101 | 21.203125)    => (001.10000 | 1.5)             
    1358 => 48,           -- (010101.001110 | 21.21875)     => (001.10000 | 1.5)             
    1359 => 48,           -- (010101.001111 | 21.234375)    => (001.10000 | 1.5)             
    1360 => 48,           -- (010101.010000 | 21.25)        => (001.10000 | 1.5)             
    1361 => 48,           -- (010101.010001 | 21.265625)    => (001.10000 | 1.5)             
    1362 => 48,           -- (010101.010010 | 21.28125)     => (001.10000 | 1.5)             
    1363 => 48,           -- (010101.010011 | 21.296875)    => (001.10000 | 1.5)             
    1364 => 48,           -- (010101.010100 | 21.3125)      => (001.10000 | 1.5)             
    1365 => 48,           -- (010101.010101 | 21.328125)    => (001.10000 | 1.5)             
    1366 => 48,           -- (010101.010110 | 21.34375)     => (001.10000 | 1.5)             
    1367 => 48,           -- (010101.010111 | 21.359375)    => (001.10000 | 1.5)             
    1368 => 48,           -- (010101.011000 | 21.375)       => (001.10000 | 1.5)             
    1369 => 48,           -- (010101.011001 | 21.390625)    => (001.10000 | 1.5)             
    1370 => 48,           -- (010101.011010 | 21.40625)     => (001.10000 | 1.5)             
    1371 => 48,           -- (010101.011011 | 21.421875)    => (001.10000 | 1.5)             
    1372 => 48,           -- (010101.011100 | 21.4375)      => (001.10000 | 1.5)             
    1373 => 48,           -- (010101.011101 | 21.453125)    => (001.10000 | 1.5)             
    1374 => 48,           -- (010101.011110 | 21.46875)     => (001.10000 | 1.5)             
    1375 => 48,           -- (010101.011111 | 21.484375)    => (001.10000 | 1.5)             
    1376 => 48,           -- (010101.100000 | 21.5)         => (001.10000 | 1.5)             
    1377 => 48,           -- (010101.100001 | 21.515625)    => (001.10000 | 1.5)             
    1378 => 48,           -- (010101.100010 | 21.53125)     => (001.10000 | 1.5)             
    1379 => 48,           -- (010101.100011 | 21.546875)    => (001.10000 | 1.5)             
    1380 => 48,           -- (010101.100100 | 21.5625)      => (001.10000 | 1.5)             
    1381 => 48,           -- (010101.100101 | 21.578125)    => (001.10000 | 1.5)             
    1382 => 48,           -- (010101.100110 | 21.59375)     => (001.10000 | 1.5)             
    1383 => 48,           -- (010101.100111 | 21.609375)    => (001.10000 | 1.5)             
    1384 => 48,           -- (010101.101000 | 21.625)       => (001.10000 | 1.5)             
    1385 => 48,           -- (010101.101001 | 21.640625)    => (001.10000 | 1.5)             
    1386 => 48,           -- (010101.101010 | 21.65625)     => (001.10000 | 1.5)             
    1387 => 48,           -- (010101.101011 | 21.671875)    => (001.10000 | 1.5)             
    1388 => 48,           -- (010101.101100 | 21.6875)      => (001.10000 | 1.5)             
    1389 => 48,           -- (010101.101101 | 21.703125)    => (001.10000 | 1.5)             
    1390 => 48,           -- (010101.101110 | 21.71875)     => (001.10000 | 1.5)             
    1391 => 48,           -- (010101.101111 | 21.734375)    => (001.10000 | 1.5)             
    1392 => 48,           -- (010101.110000 | 21.75)        => (001.10000 | 1.5)             
    1393 => 48,           -- (010101.110001 | 21.765625)    => (001.10000 | 1.5)             
    1394 => 48,           -- (010101.110010 | 21.78125)     => (001.10000 | 1.5)             
    1395 => 48,           -- (010101.110011 | 21.796875)    => (001.10000 | 1.5)             
    1396 => 48,           -- (010101.110100 | 21.8125)      => (001.10000 | 1.5)             
    1397 => 48,           -- (010101.110101 | 21.828125)    => (001.10000 | 1.5)             
    1398 => 48,           -- (010101.110110 | 21.84375)     => (001.10000 | 1.5)             
    1399 => 48,           -- (010101.110111 | 21.859375)    => (001.10000 | 1.5)             
    1400 => 48,           -- (010101.111000 | 21.875)       => (001.10000 | 1.5)             
    1401 => 48,           -- (010101.111001 | 21.890625)    => (001.10000 | 1.5)             
    1402 => 48,           -- (010101.111010 | 21.90625)     => (001.10000 | 1.5)             
    1403 => 48,           -- (010101.111011 | 21.921875)    => (001.10000 | 1.5)             
    1404 => 48,           -- (010101.111100 | 21.9375)      => (001.10000 | 1.5)             
    1405 => 48,           -- (010101.111101 | 21.953125)    => (001.10000 | 1.5)             
    1406 => 48,           -- (010101.111110 | 21.96875)     => (001.10000 | 1.5)             
    1407 => 48,           -- (010101.111111 | 21.984375)    => (001.10000 | 1.5)             
    1408 => 48,           -- (010110.000000 | 22.0)         => (001.10000 | 1.5)             
    1409 => 48,           -- (010110.000001 | 22.015625)    => (001.10000 | 1.5)             
    1410 => 48,           -- (010110.000010 | 22.03125)     => (001.10000 | 1.5)             
    1411 => 48,           -- (010110.000011 | 22.046875)    => (001.10000 | 1.5)             
    1412 => 48,           -- (010110.000100 | 22.0625)      => (001.10000 | 1.5)             
    1413 => 48,           -- (010110.000101 | 22.078125)    => (001.10000 | 1.5)             
    1414 => 48,           -- (010110.000110 | 22.09375)     => (001.10000 | 1.5)             
    1415 => 48,           -- (010110.000111 | 22.109375)    => (001.10000 | 1.5)             
    1416 => 48,           -- (010110.001000 | 22.125)       => (001.10000 | 1.5)             
    1417 => 48,           -- (010110.001001 | 22.140625)    => (001.10000 | 1.5)             
    1418 => 48,           -- (010110.001010 | 22.15625)     => (001.10000 | 1.5)             
    1419 => 48,           -- (010110.001011 | 22.171875)    => (001.10000 | 1.5)             
    1420 => 48,           -- (010110.001100 | 22.1875)      => (001.10000 | 1.5)             
    1421 => 48,           -- (010110.001101 | 22.203125)    => (001.10000 | 1.5)             
    1422 => 48,           -- (010110.001110 | 22.21875)     => (001.10000 | 1.5)             
    1423 => 48,           -- (010110.001111 | 22.234375)    => (001.10000 | 1.5)             
    1424 => 48,           -- (010110.010000 | 22.25)        => (001.10000 | 1.5)             
    1425 => 48,           -- (010110.010001 | 22.265625)    => (001.10000 | 1.5)             
    1426 => 48,           -- (010110.010010 | 22.28125)     => (001.10000 | 1.5)             
    1427 => 48,           -- (010110.010011 | 22.296875)    => (001.10000 | 1.5)             
    1428 => 48,           -- (010110.010100 | 22.3125)      => (001.10000 | 1.5)             
    1429 => 48,           -- (010110.010101 | 22.328125)    => (001.10000 | 1.5)             
    1430 => 48,           -- (010110.010110 | 22.34375)     => (001.10000 | 1.5)             
    1431 => 48,           -- (010110.010111 | 22.359375)    => (001.10000 | 1.5)             
    1432 => 48,           -- (010110.011000 | 22.375)       => (001.10000 | 1.5)             
    1433 => 48,           -- (010110.011001 | 22.390625)    => (001.10000 | 1.5)             
    1434 => 48,           -- (010110.011010 | 22.40625)     => (001.10000 | 1.5)             
    1435 => 48,           -- (010110.011011 | 22.421875)    => (001.10000 | 1.5)             
    1436 => 48,           -- (010110.011100 | 22.4375)      => (001.10000 | 1.5)             
    1437 => 48,           -- (010110.011101 | 22.453125)    => (001.10000 | 1.5)             
    1438 => 48,           -- (010110.011110 | 22.46875)     => (001.10000 | 1.5)             
    1439 => 48,           -- (010110.011111 | 22.484375)    => (001.10000 | 1.5)             
    1440 => 48,           -- (010110.100000 | 22.5)         => (001.10000 | 1.5)             
    1441 => 48,           -- (010110.100001 | 22.515625)    => (001.10000 | 1.5)             
    1442 => 48,           -- (010110.100010 | 22.53125)     => (001.10000 | 1.5)             
    1443 => 48,           -- (010110.100011 | 22.546875)    => (001.10000 | 1.5)             
    1444 => 48,           -- (010110.100100 | 22.5625)      => (001.10000 | 1.5)             
    1445 => 48,           -- (010110.100101 | 22.578125)    => (001.10000 | 1.5)             
    1446 => 48,           -- (010110.100110 | 22.59375)     => (001.10000 | 1.5)             
    1447 => 48,           -- (010110.100111 | 22.609375)    => (001.10000 | 1.5)             
    1448 => 48,           -- (010110.101000 | 22.625)       => (001.10000 | 1.5)             
    1449 => 48,           -- (010110.101001 | 22.640625)    => (001.10000 | 1.5)             
    1450 => 48,           -- (010110.101010 | 22.65625)     => (001.10000 | 1.5)             
    1451 => 48,           -- (010110.101011 | 22.671875)    => (001.10000 | 1.5)             
    1452 => 48,           -- (010110.101100 | 22.6875)      => (001.10000 | 1.5)             
    1453 => 48,           -- (010110.101101 | 22.703125)    => (001.10000 | 1.5)             
    1454 => 48,           -- (010110.101110 | 22.71875)     => (001.10000 | 1.5)             
    1455 => 48,           -- (010110.101111 | 22.734375)    => (001.10000 | 1.5)             
    1456 => 48,           -- (010110.110000 | 22.75)        => (001.10000 | 1.5)             
    1457 => 48,           -- (010110.110001 | 22.765625)    => (001.10000 | 1.5)             
    1458 => 48,           -- (010110.110010 | 22.78125)     => (001.10000 | 1.5)             
    1459 => 48,           -- (010110.110011 | 22.796875)    => (001.10000 | 1.5)             
    1460 => 48,           -- (010110.110100 | 22.8125)      => (001.10000 | 1.5)             
    1461 => 48,           -- (010110.110101 | 22.828125)    => (001.10000 | 1.5)             
    1462 => 48,           -- (010110.110110 | 22.84375)     => (001.10000 | 1.5)             
    1463 => 48,           -- (010110.110111 | 22.859375)    => (001.10000 | 1.5)             
    1464 => 48,           -- (010110.111000 | 22.875)       => (001.10000 | 1.5)             
    1465 => 48,           -- (010110.111001 | 22.890625)    => (001.10000 | 1.5)             
    1466 => 48,           -- (010110.111010 | 22.90625)     => (001.10000 | 1.5)             
    1467 => 48,           -- (010110.111011 | 22.921875)    => (001.10000 | 1.5)             
    1468 => 48,           -- (010110.111100 | 22.9375)      => (001.10000 | 1.5)             
    1469 => 48,           -- (010110.111101 | 22.953125)    => (001.10000 | 1.5)             
    1470 => 48,           -- (010110.111110 | 22.96875)     => (001.10000 | 1.5)             
    1471 => 48,           -- (010110.111111 | 22.984375)    => (001.10000 | 1.5)             
    1472 => 48,           -- (010111.000000 | 23.0)         => (001.10000 | 1.5)             
    1473 => 48,           -- (010111.000001 | 23.015625)    => (001.10000 | 1.5)             
    1474 => 48,           -- (010111.000010 | 23.03125)     => (001.10000 | 1.5)             
    1475 => 48,           -- (010111.000011 | 23.046875)    => (001.10000 | 1.5)             
    1476 => 48,           -- (010111.000100 | 23.0625)      => (001.10000 | 1.5)             
    1477 => 48,           -- (010111.000101 | 23.078125)    => (001.10000 | 1.5)             
    1478 => 48,           -- (010111.000110 | 23.09375)     => (001.10000 | 1.5)             
    1479 => 48,           -- (010111.000111 | 23.109375)    => (001.10000 | 1.5)             
    1480 => 48,           -- (010111.001000 | 23.125)       => (001.10000 | 1.5)             
    1481 => 48,           -- (010111.001001 | 23.140625)    => (001.10000 | 1.5)             
    1482 => 48,           -- (010111.001010 | 23.15625)     => (001.10000 | 1.5)             
    1483 => 48,           -- (010111.001011 | 23.171875)    => (001.10000 | 1.5)             
    1484 => 48,           -- (010111.001100 | 23.1875)      => (001.10000 | 1.5)             
    1485 => 48,           -- (010111.001101 | 23.203125)    => (001.10000 | 1.5)             
    1486 => 48,           -- (010111.001110 | 23.21875)     => (001.10000 | 1.5)             
    1487 => 48,           -- (010111.001111 | 23.234375)    => (001.10000 | 1.5)             
    1488 => 48,           -- (010111.010000 | 23.25)        => (001.10000 | 1.5)             
    1489 => 48,           -- (010111.010001 | 23.265625)    => (001.10000 | 1.5)             
    1490 => 48,           -- (010111.010010 | 23.28125)     => (001.10000 | 1.5)             
    1491 => 48,           -- (010111.010011 | 23.296875)    => (001.10000 | 1.5)             
    1492 => 48,           -- (010111.010100 | 23.3125)      => (001.10000 | 1.5)             
    1493 => 48,           -- (010111.010101 | 23.328125)    => (001.10000 | 1.5)             
    1494 => 48,           -- (010111.010110 | 23.34375)     => (001.10000 | 1.5)             
    1495 => 48,           -- (010111.010111 | 23.359375)    => (001.10000 | 1.5)             
    1496 => 48,           -- (010111.011000 | 23.375)       => (001.10000 | 1.5)             
    1497 => 48,           -- (010111.011001 | 23.390625)    => (001.10000 | 1.5)             
    1498 => 48,           -- (010111.011010 | 23.40625)     => (001.10000 | 1.5)             
    1499 => 48,           -- (010111.011011 | 23.421875)    => (001.10000 | 1.5)             
    1500 => 48,           -- (010111.011100 | 23.4375)      => (001.10000 | 1.5)             
    1501 => 48,           -- (010111.011101 | 23.453125)    => (001.10000 | 1.5)             
    1502 => 48,           -- (010111.011110 | 23.46875)     => (001.10000 | 1.5)             
    1503 => 48,           -- (010111.011111 | 23.484375)    => (001.10000 | 1.5)             
    1504 => 48,           -- (010111.100000 | 23.5)         => (001.10000 | 1.5)             
    1505 => 48,           -- (010111.100001 | 23.515625)    => (001.10000 | 1.5)             
    1506 => 48,           -- (010111.100010 | 23.53125)     => (001.10000 | 1.5)             
    1507 => 48,           -- (010111.100011 | 23.546875)    => (001.10000 | 1.5)             
    1508 => 48,           -- (010111.100100 | 23.5625)      => (001.10000 | 1.5)             
    1509 => 48,           -- (010111.100101 | 23.578125)    => (001.10000 | 1.5)             
    1510 => 48,           -- (010111.100110 | 23.59375)     => (001.10000 | 1.5)             
    1511 => 48,           -- (010111.100111 | 23.609375)    => (001.10000 | 1.5)             
    1512 => 48,           -- (010111.101000 | 23.625)       => (001.10000 | 1.5)             
    1513 => 48,           -- (010111.101001 | 23.640625)    => (001.10000 | 1.5)             
    1514 => 48,           -- (010111.101010 | 23.65625)     => (001.10000 | 1.5)             
    1515 => 48,           -- (010111.101011 | 23.671875)    => (001.10000 | 1.5)             
    1516 => 48,           -- (010111.101100 | 23.6875)      => (001.10000 | 1.5)             
    1517 => 48,           -- (010111.101101 | 23.703125)    => (001.10000 | 1.5)             
    1518 => 48,           -- (010111.101110 | 23.71875)     => (001.10000 | 1.5)             
    1519 => 48,           -- (010111.101111 | 23.734375)    => (001.10000 | 1.5)             
    1520 => 48,           -- (010111.110000 | 23.75)        => (001.10000 | 1.5)             
    1521 => 48,           -- (010111.110001 | 23.765625)    => (001.10000 | 1.5)             
    1522 => 48,           -- (010111.110010 | 23.78125)     => (001.10000 | 1.5)             
    1523 => 48,           -- (010111.110011 | 23.796875)    => (001.10000 | 1.5)             
    1524 => 48,           -- (010111.110100 | 23.8125)      => (001.10000 | 1.5)             
    1525 => 48,           -- (010111.110101 | 23.828125)    => (001.10000 | 1.5)             
    1526 => 48,           -- (010111.110110 | 23.84375)     => (001.10000 | 1.5)             
    1527 => 48,           -- (010111.110111 | 23.859375)    => (001.10000 | 1.5)             
    1528 => 48,           -- (010111.111000 | 23.875)       => (001.10000 | 1.5)             
    1529 => 48,           -- (010111.111001 | 23.890625)    => (001.10000 | 1.5)             
    1530 => 48,           -- (010111.111010 | 23.90625)     => (001.10000 | 1.5)             
    1531 => 48,           -- (010111.111011 | 23.921875)    => (001.10000 | 1.5)             
    1532 => 48,           -- (010111.111100 | 23.9375)      => (001.10000 | 1.5)             
    1533 => 48,           -- (010111.111101 | 23.953125)    => (001.10000 | 1.5)             
    1534 => 48,           -- (010111.111110 | 23.96875)     => (001.10000 | 1.5)             
    1535 => 48,           -- (010111.111111 | 23.984375)    => (001.10000 | 1.5)             
    1536 => 48,           -- (011000.000000 | 24.0)         => (001.10000 | 1.5)             
    1537 => 48,           -- (011000.000001 | 24.015625)    => (001.10000 | 1.5)             
    1538 => 48,           -- (011000.000010 | 24.03125)     => (001.10000 | 1.5)             
    1539 => 48,           -- (011000.000011 | 24.046875)    => (001.10000 | 1.5)             
    1540 => 48,           -- (011000.000100 | 24.0625)      => (001.10000 | 1.5)             
    1541 => 48,           -- (011000.000101 | 24.078125)    => (001.10000 | 1.5)             
    1542 => 48,           -- (011000.000110 | 24.09375)     => (001.10000 | 1.5)             
    1543 => 48,           -- (011000.000111 | 24.109375)    => (001.10000 | 1.5)             
    1544 => 48,           -- (011000.001000 | 24.125)       => (001.10000 | 1.5)             
    1545 => 48,           -- (011000.001001 | 24.140625)    => (001.10000 | 1.5)             
    1546 => 48,           -- (011000.001010 | 24.15625)     => (001.10000 | 1.5)             
    1547 => 48,           -- (011000.001011 | 24.171875)    => (001.10000 | 1.5)             
    1548 => 48,           -- (011000.001100 | 24.1875)      => (001.10000 | 1.5)             
    1549 => 48,           -- (011000.001101 | 24.203125)    => (001.10000 | 1.5)             
    1550 => 48,           -- (011000.001110 | 24.21875)     => (001.10000 | 1.5)             
    1551 => 48,           -- (011000.001111 | 24.234375)    => (001.10000 | 1.5)             
    1552 => 48,           -- (011000.010000 | 24.25)        => (001.10000 | 1.5)             
    1553 => 48,           -- (011000.010001 | 24.265625)    => (001.10000 | 1.5)             
    1554 => 48,           -- (011000.010010 | 24.28125)     => (001.10000 | 1.5)             
    1555 => 48,           -- (011000.010011 | 24.296875)    => (001.10000 | 1.5)             
    1556 => 48,           -- (011000.010100 | 24.3125)      => (001.10000 | 1.5)             
    1557 => 48,           -- (011000.010101 | 24.328125)    => (001.10000 | 1.5)             
    1558 => 48,           -- (011000.010110 | 24.34375)     => (001.10000 | 1.5)             
    1559 => 48,           -- (011000.010111 | 24.359375)    => (001.10000 | 1.5)             
    1560 => 48,           -- (011000.011000 | 24.375)       => (001.10000 | 1.5)             
    1561 => 48,           -- (011000.011001 | 24.390625)    => (001.10000 | 1.5)             
    1562 => 48,           -- (011000.011010 | 24.40625)     => (001.10000 | 1.5)             
    1563 => 48,           -- (011000.011011 | 24.421875)    => (001.10000 | 1.5)             
    1564 => 48,           -- (011000.011100 | 24.4375)      => (001.10000 | 1.5)             
    1565 => 48,           -- (011000.011101 | 24.453125)    => (001.10000 | 1.5)             
    1566 => 48,           -- (011000.011110 | 24.46875)     => (001.10000 | 1.5)             
    1567 => 48,           -- (011000.011111 | 24.484375)    => (001.10000 | 1.5)             
    1568 => 48,           -- (011000.100000 | 24.5)         => (001.10000 | 1.5)             
    1569 => 48,           -- (011000.100001 | 24.515625)    => (001.10000 | 1.5)             
    1570 => 48,           -- (011000.100010 | 24.53125)     => (001.10000 | 1.5)             
    1571 => 48,           -- (011000.100011 | 24.546875)    => (001.10000 | 1.5)             
    1572 => 48,           -- (011000.100100 | 24.5625)      => (001.10000 | 1.5)             
    1573 => 48,           -- (011000.100101 | 24.578125)    => (001.10000 | 1.5)             
    1574 => 48,           -- (011000.100110 | 24.59375)     => (001.10000 | 1.5)             
    1575 => 48,           -- (011000.100111 | 24.609375)    => (001.10000 | 1.5)             
    1576 => 48,           -- (011000.101000 | 24.625)       => (001.10000 | 1.5)             
    1577 => 48,           -- (011000.101001 | 24.640625)    => (001.10000 | 1.5)             
    1578 => 48,           -- (011000.101010 | 24.65625)     => (001.10000 | 1.5)             
    1579 => 48,           -- (011000.101011 | 24.671875)    => (001.10000 | 1.5)             
    1580 => 48,           -- (011000.101100 | 24.6875)      => (001.10000 | 1.5)             
    1581 => 48,           -- (011000.101101 | 24.703125)    => (001.10000 | 1.5)             
    1582 => 48,           -- (011000.101110 | 24.71875)     => (001.10000 | 1.5)             
    1583 => 48,           -- (011000.101111 | 24.734375)    => (001.10000 | 1.5)             
    1584 => 48,           -- (011000.110000 | 24.75)        => (001.10000 | 1.5)             
    1585 => 48,           -- (011000.110001 | 24.765625)    => (001.10000 | 1.5)             
    1586 => 48,           -- (011000.110010 | 24.78125)     => (001.10000 | 1.5)             
    1587 => 48,           -- (011000.110011 | 24.796875)    => (001.10000 | 1.5)             
    1588 => 48,           -- (011000.110100 | 24.8125)      => (001.10000 | 1.5)             
    1589 => 48,           -- (011000.110101 | 24.828125)    => (001.10000 | 1.5)             
    1590 => 48,           -- (011000.110110 | 24.84375)     => (001.10000 | 1.5)             
    1591 => 48,           -- (011000.110111 | 24.859375)    => (001.10000 | 1.5)             
    1592 => 48,           -- (011000.111000 | 24.875)       => (001.10000 | 1.5)             
    1593 => 48,           -- (011000.111001 | 24.890625)    => (001.10000 | 1.5)             
    1594 => 48,           -- (011000.111010 | 24.90625)     => (001.10000 | 1.5)             
    1595 => 48,           -- (011000.111011 | 24.921875)    => (001.10000 | 1.5)             
    1596 => 48,           -- (011000.111100 | 24.9375)      => (001.10000 | 1.5)             
    1597 => 48,           -- (011000.111101 | 24.953125)    => (001.10000 | 1.5)             
    1598 => 48,           -- (011000.111110 | 24.96875)     => (001.10000 | 1.5)             
    1599 => 48,           -- (011000.111111 | 24.984375)    => (001.10000 | 1.5)             
    1600 => 48,           -- (011001.000000 | 25.0)         => (001.10000 | 1.5)             
    1601 => 48,           -- (011001.000001 | 25.015625)    => (001.10000 | 1.5)             
    1602 => 48,           -- (011001.000010 | 25.03125)     => (001.10000 | 1.5)             
    1603 => 48,           -- (011001.000011 | 25.046875)    => (001.10000 | 1.5)             
    1604 => 48,           -- (011001.000100 | 25.0625)      => (001.10000 | 1.5)             
    1605 => 48,           -- (011001.000101 | 25.078125)    => (001.10000 | 1.5)             
    1606 => 48,           -- (011001.000110 | 25.09375)     => (001.10000 | 1.5)             
    1607 => 48,           -- (011001.000111 | 25.109375)    => (001.10000 | 1.5)             
    1608 => 48,           -- (011001.001000 | 25.125)       => (001.10000 | 1.5)             
    1609 => 48,           -- (011001.001001 | 25.140625)    => (001.10000 | 1.5)             
    1610 => 48,           -- (011001.001010 | 25.15625)     => (001.10000 | 1.5)             
    1611 => 48,           -- (011001.001011 | 25.171875)    => (001.10000 | 1.5)             
    1612 => 48,           -- (011001.001100 | 25.1875)      => (001.10000 | 1.5)             
    1613 => 48,           -- (011001.001101 | 25.203125)    => (001.10000 | 1.5)             
    1614 => 48,           -- (011001.001110 | 25.21875)     => (001.10000 | 1.5)             
    1615 => 48,           -- (011001.001111 | 25.234375)    => (001.10000 | 1.5)             
    1616 => 48,           -- (011001.010000 | 25.25)        => (001.10000 | 1.5)             
    1617 => 48,           -- (011001.010001 | 25.265625)    => (001.10000 | 1.5)             
    1618 => 49,           -- (011001.010010 | 25.28125)     => (001.10001 | 1.53125)         
    1619 => 49,           -- (011001.010011 | 25.296875)    => (001.10001 | 1.53125)         
    1620 => 49,           -- (011001.010100 | 25.3125)      => (001.10001 | 1.53125)         
    1621 => 49,           -- (011001.010101 | 25.328125)    => (001.10001 | 1.53125)         
    1622 => 49,           -- (011001.010110 | 25.34375)     => (001.10001 | 1.53125)         
    1623 => 49,           -- (011001.010111 | 25.359375)    => (001.10001 | 1.53125)         
    1624 => 49,           -- (011001.011000 | 25.375)       => (001.10001 | 1.53125)         
    1625 => 49,           -- (011001.011001 | 25.390625)    => (001.10001 | 1.53125)         
    1626 => 49,           -- (011001.011010 | 25.40625)     => (001.10001 | 1.53125)         
    1627 => 49,           -- (011001.011011 | 25.421875)    => (001.10001 | 1.53125)         
    1628 => 49,           -- (011001.011100 | 25.4375)      => (001.10001 | 1.53125)         
    1629 => 49,           -- (011001.011101 | 25.453125)    => (001.10001 | 1.53125)         
    1630 => 49,           -- (011001.011110 | 25.46875)     => (001.10001 | 1.53125)         
    1631 => 49,           -- (011001.011111 | 25.484375)    => (001.10001 | 1.53125)         
    1632 => 49,           -- (011001.100000 | 25.5)         => (001.10001 | 1.53125)         
    1633 => 49,           -- (011001.100001 | 25.515625)    => (001.10001 | 1.53125)         
    1634 => 49,           -- (011001.100010 | 25.53125)     => (001.10001 | 1.53125)         
    1635 => 49,           -- (011001.100011 | 25.546875)    => (001.10001 | 1.53125)         
    1636 => 49,           -- (011001.100100 | 25.5625)      => (001.10001 | 1.53125)         
    1637 => 49,           -- (011001.100101 | 25.578125)    => (001.10001 | 1.53125)         
    1638 => 49,           -- (011001.100110 | 25.59375)     => (001.10001 | 1.53125)         
    1639 => 49,           -- (011001.100111 | 25.609375)    => (001.10001 | 1.53125)         
    1640 => 49,           -- (011001.101000 | 25.625)       => (001.10001 | 1.53125)         
    1641 => 49,           -- (011001.101001 | 25.640625)    => (001.10001 | 1.53125)         
    1642 => 49,           -- (011001.101010 | 25.65625)     => (001.10001 | 1.53125)         
    1643 => 49,           -- (011001.101011 | 25.671875)    => (001.10001 | 1.53125)         
    1644 => 49,           -- (011001.101100 | 25.6875)      => (001.10001 | 1.53125)         
    1645 => 49,           -- (011001.101101 | 25.703125)    => (001.10001 | 1.53125)         
    1646 => 49,           -- (011001.101110 | 25.71875)     => (001.10001 | 1.53125)         
    1647 => 49,           -- (011001.101111 | 25.734375)    => (001.10001 | 1.53125)         
    1648 => 49,           -- (011001.110000 | 25.75)        => (001.10001 | 1.53125)         
    1649 => 49,           -- (011001.110001 | 25.765625)    => (001.10001 | 1.53125)         
    1650 => 49,           -- (011001.110010 | 25.78125)     => (001.10001 | 1.53125)         
    1651 => 49,           -- (011001.110011 | 25.796875)    => (001.10001 | 1.53125)         
    1652 => 49,           -- (011001.110100 | 25.8125)      => (001.10001 | 1.53125)         
    1653 => 49,           -- (011001.110101 | 25.828125)    => (001.10001 | 1.53125)         
    1654 => 49,           -- (011001.110110 | 25.84375)     => (001.10001 | 1.53125)         
    1655 => 49,           -- (011001.110111 | 25.859375)    => (001.10001 | 1.53125)         
    1656 => 49,           -- (011001.111000 | 25.875)       => (001.10001 | 1.53125)         
    1657 => 49,           -- (011001.111001 | 25.890625)    => (001.10001 | 1.53125)         
    1658 => 49,           -- (011001.111010 | 25.90625)     => (001.10001 | 1.53125)         
    1659 => 49,           -- (011001.111011 | 25.921875)    => (001.10001 | 1.53125)         
    1660 => 49,           -- (011001.111100 | 25.9375)      => (001.10001 | 1.53125)         
    1661 => 49,           -- (011001.111101 | 25.953125)    => (001.10001 | 1.53125)         
    1662 => 49,           -- (011001.111110 | 25.96875)     => (001.10001 | 1.53125)         
    1663 => 49,           -- (011001.111111 | 25.984375)    => (001.10001 | 1.53125)         
    1664 => 49,           -- (011010.000000 | 26.0)         => (001.10001 | 1.53125)         
    1665 => 49,           -- (011010.000001 | 26.015625)    => (001.10001 | 1.53125)         
    1666 => 49,           -- (011010.000010 | 26.03125)     => (001.10001 | 1.53125)         
    1667 => 49,           -- (011010.000011 | 26.046875)    => (001.10001 | 1.53125)         
    1668 => 49,           -- (011010.000100 | 26.0625)      => (001.10001 | 1.53125)         
    1669 => 49,           -- (011010.000101 | 26.078125)    => (001.10001 | 1.53125)         
    1670 => 49,           -- (011010.000110 | 26.09375)     => (001.10001 | 1.53125)         
    1671 => 49,           -- (011010.000111 | 26.109375)    => (001.10001 | 1.53125)         
    1672 => 49,           -- (011010.001000 | 26.125)       => (001.10001 | 1.53125)         
    1673 => 49,           -- (011010.001001 | 26.140625)    => (001.10001 | 1.53125)         
    1674 => 49,           -- (011010.001010 | 26.15625)     => (001.10001 | 1.53125)         
    1675 => 49,           -- (011010.001011 | 26.171875)    => (001.10001 | 1.53125)         
    1676 => 49,           -- (011010.001100 | 26.1875)      => (001.10001 | 1.53125)         
    1677 => 49,           -- (011010.001101 | 26.203125)    => (001.10001 | 1.53125)         
    1678 => 49,           -- (011010.001110 | 26.21875)     => (001.10001 | 1.53125)         
    1679 => 49,           -- (011010.001111 | 26.234375)    => (001.10001 | 1.53125)         
    1680 => 49,           -- (011010.010000 | 26.25)        => (001.10001 | 1.53125)         
    1681 => 49,           -- (011010.010001 | 26.265625)    => (001.10001 | 1.53125)         
    1682 => 49,           -- (011010.010010 | 26.28125)     => (001.10001 | 1.53125)         
    1683 => 49,           -- (011010.010011 | 26.296875)    => (001.10001 | 1.53125)         
    1684 => 49,           -- (011010.010100 | 26.3125)      => (001.10001 | 1.53125)         
    1685 => 49,           -- (011010.010101 | 26.328125)    => (001.10001 | 1.53125)         
    1686 => 49,           -- (011010.010110 | 26.34375)     => (001.10001 | 1.53125)         
    1687 => 49,           -- (011010.010111 | 26.359375)    => (001.10001 | 1.53125)         
    1688 => 49,           -- (011010.011000 | 26.375)       => (001.10001 | 1.53125)         
    1689 => 49,           -- (011010.011001 | 26.390625)    => (001.10001 | 1.53125)         
    1690 => 49,           -- (011010.011010 | 26.40625)     => (001.10001 | 1.53125)         
    1691 => 49,           -- (011010.011011 | 26.421875)    => (001.10001 | 1.53125)         
    1692 => 49,           -- (011010.011100 | 26.4375)      => (001.10001 | 1.53125)         
    1693 => 49,           -- (011010.011101 | 26.453125)    => (001.10001 | 1.53125)         
    1694 => 49,           -- (011010.011110 | 26.46875)     => (001.10001 | 1.53125)         
    1695 => 49,           -- (011010.011111 | 26.484375)    => (001.10001 | 1.53125)         
    1696 => 49,           -- (011010.100000 | 26.5)         => (001.10001 | 1.53125)         
    1697 => 49,           -- (011010.100001 | 26.515625)    => (001.10001 | 1.53125)         
    1698 => 49,           -- (011010.100010 | 26.53125)     => (001.10001 | 1.53125)         
    1699 => 49,           -- (011010.100011 | 26.546875)    => (001.10001 | 1.53125)         
    1700 => 49,           -- (011010.100100 | 26.5625)      => (001.10001 | 1.53125)         
    1701 => 49,           -- (011010.100101 | 26.578125)    => (001.10001 | 1.53125)         
    1702 => 49,           -- (011010.100110 | 26.59375)     => (001.10001 | 1.53125)         
    1703 => 49,           -- (011010.100111 | 26.609375)    => (001.10001 | 1.53125)         
    1704 => 49,           -- (011010.101000 | 26.625)       => (001.10001 | 1.53125)         
    1705 => 49,           -- (011010.101001 | 26.640625)    => (001.10001 | 1.53125)         
    1706 => 49,           -- (011010.101010 | 26.65625)     => (001.10001 | 1.53125)         
    1707 => 49,           -- (011010.101011 | 26.671875)    => (001.10001 | 1.53125)         
    1708 => 49,           -- (011010.101100 | 26.6875)      => (001.10001 | 1.53125)         
    1709 => 49,           -- (011010.101101 | 26.703125)    => (001.10001 | 1.53125)         
    1710 => 49,           -- (011010.101110 | 26.71875)     => (001.10001 | 1.53125)         
    1711 => 49,           -- (011010.101111 | 26.734375)    => (001.10001 | 1.53125)         
    1712 => 49,           -- (011010.110000 | 26.75)        => (001.10001 | 1.53125)         
    1713 => 49,           -- (011010.110001 | 26.765625)    => (001.10001 | 1.53125)         
    1714 => 49,           -- (011010.110010 | 26.78125)     => (001.10001 | 1.53125)         
    1715 => 49,           -- (011010.110011 | 26.796875)    => (001.10001 | 1.53125)         
    1716 => 49,           -- (011010.110100 | 26.8125)      => (001.10001 | 1.53125)         
    1717 => 49,           -- (011010.110101 | 26.828125)    => (001.10001 | 1.53125)         
    1718 => 49,           -- (011010.110110 | 26.84375)     => (001.10001 | 1.53125)         
    1719 => 49,           -- (011010.110111 | 26.859375)    => (001.10001 | 1.53125)         
    1720 => 49,           -- (011010.111000 | 26.875)       => (001.10001 | 1.53125)         
    1721 => 49,           -- (011010.111001 | 26.890625)    => (001.10001 | 1.53125)         
    1722 => 49,           -- (011010.111010 | 26.90625)     => (001.10001 | 1.53125)         
    1723 => 49,           -- (011010.111011 | 26.921875)    => (001.10001 | 1.53125)         
    1724 => 49,           -- (011010.111100 | 26.9375)      => (001.10001 | 1.53125)         
    1725 => 49,           -- (011010.111101 | 26.953125)    => (001.10001 | 1.53125)         
    1726 => 49,           -- (011010.111110 | 26.96875)     => (001.10001 | 1.53125)         
    1727 => 49,           -- (011010.111111 | 26.984375)    => (001.10001 | 1.53125)         
    1728 => 49,           -- (011011.000000 | 27.0)         => (001.10001 | 1.53125)         
    1729 => 49,           -- (011011.000001 | 27.015625)    => (001.10001 | 1.53125)         
    1730 => 49,           -- (011011.000010 | 27.03125)     => (001.10001 | 1.53125)         
    1731 => 49,           -- (011011.000011 | 27.046875)    => (001.10001 | 1.53125)         
    1732 => 49,           -- (011011.000100 | 27.0625)      => (001.10001 | 1.53125)         
    1733 => 49,           -- (011011.000101 | 27.078125)    => (001.10001 | 1.53125)         
    1734 => 49,           -- (011011.000110 | 27.09375)     => (001.10001 | 1.53125)         
    1735 => 49,           -- (011011.000111 | 27.109375)    => (001.10001 | 1.53125)         
    1736 => 49,           -- (011011.001000 | 27.125)       => (001.10001 | 1.53125)         
    1737 => 49,           -- (011011.001001 | 27.140625)    => (001.10001 | 1.53125)         
    1738 => 49,           -- (011011.001010 | 27.15625)     => (001.10001 | 1.53125)         
    1739 => 49,           -- (011011.001011 | 27.171875)    => (001.10001 | 1.53125)         
    1740 => 49,           -- (011011.001100 | 27.1875)      => (001.10001 | 1.53125)         
    1741 => 49,           -- (011011.001101 | 27.203125)    => (001.10001 | 1.53125)         
    1742 => 49,           -- (011011.001110 | 27.21875)     => (001.10001 | 1.53125)         
    1743 => 49,           -- (011011.001111 | 27.234375)    => (001.10001 | 1.53125)         
    1744 => 49,           -- (011011.010000 | 27.25)        => (001.10001 | 1.53125)         
    1745 => 49,           -- (011011.010001 | 27.265625)    => (001.10001 | 1.53125)         
    1746 => 49,           -- (011011.010010 | 27.28125)     => (001.10001 | 1.53125)         
    1747 => 49,           -- (011011.010011 | 27.296875)    => (001.10001 | 1.53125)         
    1748 => 49,           -- (011011.010100 | 27.3125)      => (001.10001 | 1.53125)         
    1749 => 49,           -- (011011.010101 | 27.328125)    => (001.10001 | 1.53125)         
    1750 => 49,           -- (011011.010110 | 27.34375)     => (001.10001 | 1.53125)         
    1751 => 49,           -- (011011.010111 | 27.359375)    => (001.10001 | 1.53125)         
    1752 => 49,           -- (011011.011000 | 27.375)       => (001.10001 | 1.53125)         
    1753 => 49,           -- (011011.011001 | 27.390625)    => (001.10001 | 1.53125)         
    1754 => 49,           -- (011011.011010 | 27.40625)     => (001.10001 | 1.53125)         
    1755 => 49,           -- (011011.011011 | 27.421875)    => (001.10001 | 1.53125)         
    1756 => 49,           -- (011011.011100 | 27.4375)      => (001.10001 | 1.53125)         
    1757 => 49,           -- (011011.011101 | 27.453125)    => (001.10001 | 1.53125)         
    1758 => 49,           -- (011011.011110 | 27.46875)     => (001.10001 | 1.53125)         
    1759 => 49,           -- (011011.011111 | 27.484375)    => (001.10001 | 1.53125)         
    1760 => 49,           -- (011011.100000 | 27.5)         => (001.10001 | 1.53125)         
    1761 => 49,           -- (011011.100001 | 27.515625)    => (001.10001 | 1.53125)         
    1762 => 49,           -- (011011.100010 | 27.53125)     => (001.10001 | 1.53125)         
    1763 => 49,           -- (011011.100011 | 27.546875)    => (001.10001 | 1.53125)         
    1764 => 49,           -- (011011.100100 | 27.5625)      => (001.10001 | 1.53125)         
    1765 => 49,           -- (011011.100101 | 27.578125)    => (001.10001 | 1.53125)         
    1766 => 49,           -- (011011.100110 | 27.59375)     => (001.10001 | 1.53125)         
    1767 => 49,           -- (011011.100111 | 27.609375)    => (001.10001 | 1.53125)         
    1768 => 49,           -- (011011.101000 | 27.625)       => (001.10001 | 1.53125)         
    1769 => 49,           -- (011011.101001 | 27.640625)    => (001.10001 | 1.53125)         
    1770 => 49,           -- (011011.101010 | 27.65625)     => (001.10001 | 1.53125)         
    1771 => 49,           -- (011011.101011 | 27.671875)    => (001.10001 | 1.53125)         
    1772 => 49,           -- (011011.101100 | 27.6875)      => (001.10001 | 1.53125)         
    1773 => 49,           -- (011011.101101 | 27.703125)    => (001.10001 | 1.53125)         
    1774 => 49,           -- (011011.101110 | 27.71875)     => (001.10001 | 1.53125)         
    1775 => 49,           -- (011011.101111 | 27.734375)    => (001.10001 | 1.53125)         
    1776 => 49,           -- (011011.110000 | 27.75)        => (001.10001 | 1.53125)         
    1777 => 49,           -- (011011.110001 | 27.765625)    => (001.10001 | 1.53125)         
    1778 => 49,           -- (011011.110010 | 27.78125)     => (001.10001 | 1.53125)         
    1779 => 49,           -- (011011.110011 | 27.796875)    => (001.10001 | 1.53125)         
    1780 => 49,           -- (011011.110100 | 27.8125)      => (001.10001 | 1.53125)         
    1781 => 49,           -- (011011.110101 | 27.828125)    => (001.10001 | 1.53125)         
    1782 => 49,           -- (011011.110110 | 27.84375)     => (001.10001 | 1.53125)         
    1783 => 49,           -- (011011.110111 | 27.859375)    => (001.10001 | 1.53125)         
    1784 => 49,           -- (011011.111000 | 27.875)       => (001.10001 | 1.53125)         
    1785 => 49,           -- (011011.111001 | 27.890625)    => (001.10001 | 1.53125)         
    1786 => 49,           -- (011011.111010 | 27.90625)     => (001.10001 | 1.53125)         
    1787 => 49,           -- (011011.111011 | 27.921875)    => (001.10001 | 1.53125)         
    1788 => 49,           -- (011011.111100 | 27.9375)      => (001.10001 | 1.53125)         
    1789 => 49,           -- (011011.111101 | 27.953125)    => (001.10001 | 1.53125)         
    1790 => 49,           -- (011011.111110 | 27.96875)     => (001.10001 | 1.53125)         
    1791 => 49,           -- (011011.111111 | 27.984375)    => (001.10001 | 1.53125)         
    1792 => 49,           -- (011100.000000 | 28.0)         => (001.10001 | 1.53125)         
    1793 => 49,           -- (011100.000001 | 28.015625)    => (001.10001 | 1.53125)         
    1794 => 49,           -- (011100.000010 | 28.03125)     => (001.10001 | 1.53125)         
    1795 => 49,           -- (011100.000011 | 28.046875)    => (001.10001 | 1.53125)         
    1796 => 49,           -- (011100.000100 | 28.0625)      => (001.10001 | 1.53125)         
    1797 => 49,           -- (011100.000101 | 28.078125)    => (001.10001 | 1.53125)         
    1798 => 49,           -- (011100.000110 | 28.09375)     => (001.10001 | 1.53125)         
    1799 => 49,           -- (011100.000111 | 28.109375)    => (001.10001 | 1.53125)         
    1800 => 49,           -- (011100.001000 | 28.125)       => (001.10001 | 1.53125)         
    1801 => 49,           -- (011100.001001 | 28.140625)    => (001.10001 | 1.53125)         
    1802 => 49,           -- (011100.001010 | 28.15625)     => (001.10001 | 1.53125)         
    1803 => 49,           -- (011100.001011 | 28.171875)    => (001.10001 | 1.53125)         
    1804 => 49,           -- (011100.001100 | 28.1875)      => (001.10001 | 1.53125)         
    1805 => 49,           -- (011100.001101 | 28.203125)    => (001.10001 | 1.53125)         
    1806 => 49,           -- (011100.001110 | 28.21875)     => (001.10001 | 1.53125)         
    1807 => 49,           -- (011100.001111 | 28.234375)    => (001.10001 | 1.53125)         
    1808 => 49,           -- (011100.010000 | 28.25)        => (001.10001 | 1.53125)         
    1809 => 49,           -- (011100.010001 | 28.265625)    => (001.10001 | 1.53125)         
    1810 => 49,           -- (011100.010010 | 28.28125)     => (001.10001 | 1.53125)         
    1811 => 49,           -- (011100.010011 | 28.296875)    => (001.10001 | 1.53125)         
    1812 => 49,           -- (011100.010100 | 28.3125)      => (001.10001 | 1.53125)         
    1813 => 49,           -- (011100.010101 | 28.328125)    => (001.10001 | 1.53125)         
    1814 => 49,           -- (011100.010110 | 28.34375)     => (001.10001 | 1.53125)         
    1815 => 49,           -- (011100.010111 | 28.359375)    => (001.10001 | 1.53125)         
    1816 => 49,           -- (011100.011000 | 28.375)       => (001.10001 | 1.53125)         
    1817 => 49,           -- (011100.011001 | 28.390625)    => (001.10001 | 1.53125)         
    1818 => 49,           -- (011100.011010 | 28.40625)     => (001.10001 | 1.53125)         
    1819 => 49,           -- (011100.011011 | 28.421875)    => (001.10001 | 1.53125)         
    1820 => 49,           -- (011100.011100 | 28.4375)      => (001.10001 | 1.53125)         
    1821 => 49,           -- (011100.011101 | 28.453125)    => (001.10001 | 1.53125)         
    1822 => 49,           -- (011100.011110 | 28.46875)     => (001.10001 | 1.53125)         
    1823 => 49,           -- (011100.011111 | 28.484375)    => (001.10001 | 1.53125)         
    1824 => 49,           -- (011100.100000 | 28.5)         => (001.10001 | 1.53125)         
    1825 => 49,           -- (011100.100001 | 28.515625)    => (001.10001 | 1.53125)         
    1826 => 49,           -- (011100.100010 | 28.53125)     => (001.10001 | 1.53125)         
    1827 => 49,           -- (011100.100011 | 28.546875)    => (001.10001 | 1.53125)         
    1828 => 49,           -- (011100.100100 | 28.5625)      => (001.10001 | 1.53125)         
    1829 => 49,           -- (011100.100101 | 28.578125)    => (001.10001 | 1.53125)         
    1830 => 49,           -- (011100.100110 | 28.59375)     => (001.10001 | 1.53125)         
    1831 => 49,           -- (011100.100111 | 28.609375)    => (001.10001 | 1.53125)         
    1832 => 49,           -- (011100.101000 | 28.625)       => (001.10001 | 1.53125)         
    1833 => 49,           -- (011100.101001 | 28.640625)    => (001.10001 | 1.53125)         
    1834 => 49,           -- (011100.101010 | 28.65625)     => (001.10001 | 1.53125)         
    1835 => 49,           -- (011100.101011 | 28.671875)    => (001.10001 | 1.53125)         
    1836 => 49,           -- (011100.101100 | 28.6875)      => (001.10001 | 1.53125)         
    1837 => 49,           -- (011100.101101 | 28.703125)    => (001.10001 | 1.53125)         
    1838 => 49,           -- (011100.101110 | 28.71875)     => (001.10001 | 1.53125)         
    1839 => 49,           -- (011100.101111 | 28.734375)    => (001.10001 | 1.53125)         
    1840 => 49,           -- (011100.110000 | 28.75)        => (001.10001 | 1.53125)         
    1841 => 49,           -- (011100.110001 | 28.765625)    => (001.10001 | 1.53125)         
    1842 => 49,           -- (011100.110010 | 28.78125)     => (001.10001 | 1.53125)         
    1843 => 49,           -- (011100.110011 | 28.796875)    => (001.10001 | 1.53125)         
    1844 => 49,           -- (011100.110100 | 28.8125)      => (001.10001 | 1.53125)         
    1845 => 49,           -- (011100.110101 | 28.828125)    => (001.10001 | 1.53125)         
    1846 => 49,           -- (011100.110110 | 28.84375)     => (001.10001 | 1.53125)         
    1847 => 49,           -- (011100.110111 | 28.859375)    => (001.10001 | 1.53125)         
    1848 => 49,           -- (011100.111000 | 28.875)       => (001.10001 | 1.53125)         
    1849 => 49,           -- (011100.111001 | 28.890625)    => (001.10001 | 1.53125)         
    1850 => 49,           -- (011100.111010 | 28.90625)     => (001.10001 | 1.53125)         
    1851 => 49,           -- (011100.111011 | 28.921875)    => (001.10001 | 1.53125)         
    1852 => 49,           -- (011100.111100 | 28.9375)      => (001.10001 | 1.53125)         
    1853 => 49,           -- (011100.111101 | 28.953125)    => (001.10001 | 1.53125)         
    1854 => 49,           -- (011100.111110 | 28.96875)     => (001.10001 | 1.53125)         
    1855 => 49,           -- (011100.111111 | 28.984375)    => (001.10001 | 1.53125)         
    1856 => 49,           -- (011101.000000 | 29.0)         => (001.10001 | 1.53125)         
    1857 => 49,           -- (011101.000001 | 29.015625)    => (001.10001 | 1.53125)         
    1858 => 49,           -- (011101.000010 | 29.03125)     => (001.10001 | 1.53125)         
    1859 => 49,           -- (011101.000011 | 29.046875)    => (001.10001 | 1.53125)         
    1860 => 49,           -- (011101.000100 | 29.0625)      => (001.10001 | 1.53125)         
    1861 => 49,           -- (011101.000101 | 29.078125)    => (001.10001 | 1.53125)         
    1862 => 49,           -- (011101.000110 | 29.09375)     => (001.10001 | 1.53125)         
    1863 => 49,           -- (011101.000111 | 29.109375)    => (001.10001 | 1.53125)         
    1864 => 49,           -- (011101.001000 | 29.125)       => (001.10001 | 1.53125)         
    1865 => 49,           -- (011101.001001 | 29.140625)    => (001.10001 | 1.53125)         
    1866 => 49,           -- (011101.001010 | 29.15625)     => (001.10001 | 1.53125)         
    1867 => 49,           -- (011101.001011 | 29.171875)    => (001.10001 | 1.53125)         
    1868 => 49,           -- (011101.001100 | 29.1875)      => (001.10001 | 1.53125)         
    1869 => 49,           -- (011101.001101 | 29.203125)    => (001.10001 | 1.53125)         
    1870 => 49,           -- (011101.001110 | 29.21875)     => (001.10001 | 1.53125)         
    1871 => 49,           -- (011101.001111 | 29.234375)    => (001.10001 | 1.53125)         
    1872 => 49,           -- (011101.010000 | 29.25)        => (001.10001 | 1.53125)         
    1873 => 49,           -- (011101.010001 | 29.265625)    => (001.10001 | 1.53125)         
    1874 => 49,           -- (011101.010010 | 29.28125)     => (001.10001 | 1.53125)         
    1875 => 49,           -- (011101.010011 | 29.296875)    => (001.10001 | 1.53125)         
    1876 => 49,           -- (011101.010100 | 29.3125)      => (001.10001 | 1.53125)         
    1877 => 49,           -- (011101.010101 | 29.328125)    => (001.10001 | 1.53125)         
    1878 => 49,           -- (011101.010110 | 29.34375)     => (001.10001 | 1.53125)         
    1879 => 49,           -- (011101.010111 | 29.359375)    => (001.10001 | 1.53125)         
    1880 => 49,           -- (011101.011000 | 29.375)       => (001.10001 | 1.53125)         
    1881 => 49,           -- (011101.011001 | 29.390625)    => (001.10001 | 1.53125)         
    1882 => 49,           -- (011101.011010 | 29.40625)     => (001.10001 | 1.53125)         
    1883 => 49,           -- (011101.011011 | 29.421875)    => (001.10001 | 1.53125)         
    1884 => 49,           -- (011101.011100 | 29.4375)      => (001.10001 | 1.53125)         
    1885 => 49,           -- (011101.011101 | 29.453125)    => (001.10001 | 1.53125)         
    1886 => 49,           -- (011101.011110 | 29.46875)     => (001.10001 | 1.53125)         
    1887 => 49,           -- (011101.011111 | 29.484375)    => (001.10001 | 1.53125)         
    1888 => 49,           -- (011101.100000 | 29.5)         => (001.10001 | 1.53125)         
    1889 => 49,           -- (011101.100001 | 29.515625)    => (001.10001 | 1.53125)         
    1890 => 49,           -- (011101.100010 | 29.53125)     => (001.10001 | 1.53125)         
    1891 => 49,           -- (011101.100011 | 29.546875)    => (001.10001 | 1.53125)         
    1892 => 49,           -- (011101.100100 | 29.5625)      => (001.10001 | 1.53125)         
    1893 => 49,           -- (011101.100101 | 29.578125)    => (001.10001 | 1.53125)         
    1894 => 49,           -- (011101.100110 | 29.59375)     => (001.10001 | 1.53125)         
    1895 => 49,           -- (011101.100111 | 29.609375)    => (001.10001 | 1.53125)         
    1896 => 49,           -- (011101.101000 | 29.625)       => (001.10001 | 1.53125)         
    1897 => 49,           -- (011101.101001 | 29.640625)    => (001.10001 | 1.53125)         
    1898 => 49,           -- (011101.101010 | 29.65625)     => (001.10001 | 1.53125)         
    1899 => 49,           -- (011101.101011 | 29.671875)    => (001.10001 | 1.53125)         
    1900 => 49,           -- (011101.101100 | 29.6875)      => (001.10001 | 1.53125)         
    1901 => 49,           -- (011101.101101 | 29.703125)    => (001.10001 | 1.53125)         
    1902 => 49,           -- (011101.101110 | 29.71875)     => (001.10001 | 1.53125)         
    1903 => 49,           -- (011101.101111 | 29.734375)    => (001.10001 | 1.53125)         
    1904 => 49,           -- (011101.110000 | 29.75)        => (001.10001 | 1.53125)         
    1905 => 49,           -- (011101.110001 | 29.765625)    => (001.10001 | 1.53125)         
    1906 => 49,           -- (011101.110010 | 29.78125)     => (001.10001 | 1.53125)         
    1907 => 49,           -- (011101.110011 | 29.796875)    => (001.10001 | 1.53125)         
    1908 => 49,           -- (011101.110100 | 29.8125)      => (001.10001 | 1.53125)         
    1909 => 49,           -- (011101.110101 | 29.828125)    => (001.10001 | 1.53125)         
    1910 => 49,           -- (011101.110110 | 29.84375)     => (001.10001 | 1.53125)         
    1911 => 49,           -- (011101.110111 | 29.859375)    => (001.10001 | 1.53125)         
    1912 => 49,           -- (011101.111000 | 29.875)       => (001.10001 | 1.53125)         
    1913 => 49,           -- (011101.111001 | 29.890625)    => (001.10001 | 1.53125)         
    1914 => 49,           -- (011101.111010 | 29.90625)     => (001.10001 | 1.53125)         
    1915 => 49,           -- (011101.111011 | 29.921875)    => (001.10001 | 1.53125)         
    1916 => 49,           -- (011101.111100 | 29.9375)      => (001.10001 | 1.53125)         
    1917 => 49,           -- (011101.111101 | 29.953125)    => (001.10001 | 1.53125)         
    1918 => 49,           -- (011101.111110 | 29.96875)     => (001.10001 | 1.53125)         
    1919 => 49,           -- (011101.111111 | 29.984375)    => (001.10001 | 1.53125)         
    1920 => 49,           -- (011110.000000 | 30.0)         => (001.10001 | 1.53125)         
    1921 => 49,           -- (011110.000001 | 30.015625)    => (001.10001 | 1.53125)         
    1922 => 49,           -- (011110.000010 | 30.03125)     => (001.10001 | 1.53125)         
    1923 => 49,           -- (011110.000011 | 30.046875)    => (001.10001 | 1.53125)         
    1924 => 49,           -- (011110.000100 | 30.0625)      => (001.10001 | 1.53125)         
    1925 => 49,           -- (011110.000101 | 30.078125)    => (001.10001 | 1.53125)         
    1926 => 49,           -- (011110.000110 | 30.09375)     => (001.10001 | 1.53125)         
    1927 => 49,           -- (011110.000111 | 30.109375)    => (001.10001 | 1.53125)         
    1928 => 49,           -- (011110.001000 | 30.125)       => (001.10001 | 1.53125)         
    1929 => 49,           -- (011110.001001 | 30.140625)    => (001.10001 | 1.53125)         
    1930 => 49,           -- (011110.001010 | 30.15625)     => (001.10001 | 1.53125)         
    1931 => 49,           -- (011110.001011 | 30.171875)    => (001.10001 | 1.53125)         
    1932 => 49,           -- (011110.001100 | 30.1875)      => (001.10001 | 1.53125)         
    1933 => 49,           -- (011110.001101 | 30.203125)    => (001.10001 | 1.53125)         
    1934 => 49,           -- (011110.001110 | 30.21875)     => (001.10001 | 1.53125)         
    1935 => 49,           -- (011110.001111 | 30.234375)    => (001.10001 | 1.53125)         
    1936 => 49,           -- (011110.010000 | 30.25)        => (001.10001 | 1.53125)         
    1937 => 49,           -- (011110.010001 | 30.265625)    => (001.10001 | 1.53125)         
    1938 => 49,           -- (011110.010010 | 30.28125)     => (001.10001 | 1.53125)         
    1939 => 49,           -- (011110.010011 | 30.296875)    => (001.10001 | 1.53125)         
    1940 => 49,           -- (011110.010100 | 30.3125)      => (001.10001 | 1.53125)         
    1941 => 49,           -- (011110.010101 | 30.328125)    => (001.10001 | 1.53125)         
    1942 => 49,           -- (011110.010110 | 30.34375)     => (001.10001 | 1.53125)         
    1943 => 49,           -- (011110.010111 | 30.359375)    => (001.10001 | 1.53125)         
    1944 => 49,           -- (011110.011000 | 30.375)       => (001.10001 | 1.53125)         
    1945 => 49,           -- (011110.011001 | 30.390625)    => (001.10001 | 1.53125)         
    1946 => 49,           -- (011110.011010 | 30.40625)     => (001.10001 | 1.53125)         
    1947 => 49,           -- (011110.011011 | 30.421875)    => (001.10001 | 1.53125)         
    1948 => 49,           -- (011110.011100 | 30.4375)      => (001.10001 | 1.53125)         
    1949 => 49,           -- (011110.011101 | 30.453125)    => (001.10001 | 1.53125)         
    1950 => 49,           -- (011110.011110 | 30.46875)     => (001.10001 | 1.53125)         
    1951 => 49,           -- (011110.011111 | 30.484375)    => (001.10001 | 1.53125)         
    1952 => 49,           -- (011110.100000 | 30.5)         => (001.10001 | 1.53125)         
    1953 => 49,           -- (011110.100001 | 30.515625)    => (001.10001 | 1.53125)         
    1954 => 49,           -- (011110.100010 | 30.53125)     => (001.10001 | 1.53125)         
    1955 => 49,           -- (011110.100011 | 30.546875)    => (001.10001 | 1.53125)         
    1956 => 49,           -- (011110.100100 | 30.5625)      => (001.10001 | 1.53125)         
    1957 => 49,           -- (011110.100101 | 30.578125)    => (001.10001 | 1.53125)         
    1958 => 49,           -- (011110.100110 | 30.59375)     => (001.10001 | 1.53125)         
    1959 => 49,           -- (011110.100111 | 30.609375)    => (001.10001 | 1.53125)         
    1960 => 49,           -- (011110.101000 | 30.625)       => (001.10001 | 1.53125)         
    1961 => 49,           -- (011110.101001 | 30.640625)    => (001.10001 | 1.53125)         
    1962 => 49,           -- (011110.101010 | 30.65625)     => (001.10001 | 1.53125)         
    1963 => 49,           -- (011110.101011 | 30.671875)    => (001.10001 | 1.53125)         
    1964 => 49,           -- (011110.101100 | 30.6875)      => (001.10001 | 1.53125)         
    1965 => 49,           -- (011110.101101 | 30.703125)    => (001.10001 | 1.53125)         
    1966 => 49,           -- (011110.101110 | 30.71875)     => (001.10001 | 1.53125)         
    1967 => 49,           -- (011110.101111 | 30.734375)    => (001.10001 | 1.53125)         
    1968 => 49,           -- (011110.110000 | 30.75)        => (001.10001 | 1.53125)         
    1969 => 49,           -- (011110.110001 | 30.765625)    => (001.10001 | 1.53125)         
    1970 => 49,           -- (011110.110010 | 30.78125)     => (001.10001 | 1.53125)         
    1971 => 49,           -- (011110.110011 | 30.796875)    => (001.10001 | 1.53125)         
    1972 => 49,           -- (011110.110100 | 30.8125)      => (001.10001 | 1.53125)         
    1973 => 49,           -- (011110.110101 | 30.828125)    => (001.10001 | 1.53125)         
    1974 => 49,           -- (011110.110110 | 30.84375)     => (001.10001 | 1.53125)         
    1975 => 49,           -- (011110.110111 | 30.859375)    => (001.10001 | 1.53125)         
    1976 => 49,           -- (011110.111000 | 30.875)       => (001.10001 | 1.53125)         
    1977 => 49,           -- (011110.111001 | 30.890625)    => (001.10001 | 1.53125)         
    1978 => 49,           -- (011110.111010 | 30.90625)     => (001.10001 | 1.53125)         
    1979 => 49,           -- (011110.111011 | 30.921875)    => (001.10001 | 1.53125)         
    1980 => 49,           -- (011110.111100 | 30.9375)      => (001.10001 | 1.53125)         
    1981 => 49,           -- (011110.111101 | 30.953125)    => (001.10001 | 1.53125)         
    1982 => 49,           -- (011110.111110 | 30.96875)     => (001.10001 | 1.53125)         
    1983 => 49,           -- (011110.111111 | 30.984375)    => (001.10001 | 1.53125)         
    1984 => 49,           -- (011111.000000 | 31.0)         => (001.10001 | 1.53125)         
    1985 => 49,           -- (011111.000001 | 31.015625)    => (001.10001 | 1.53125)         
    1986 => 49,           -- (011111.000010 | 31.03125)     => (001.10001 | 1.53125)         
    1987 => 49,           -- (011111.000011 | 31.046875)    => (001.10001 | 1.53125)         
    1988 => 49,           -- (011111.000100 | 31.0625)      => (001.10001 | 1.53125)         
    1989 => 49,           -- (011111.000101 | 31.078125)    => (001.10001 | 1.53125)         
    1990 => 49,           -- (011111.000110 | 31.09375)     => (001.10001 | 1.53125)         
    1991 => 49,           -- (011111.000111 | 31.109375)    => (001.10001 | 1.53125)         
    1992 => 49,           -- (011111.001000 | 31.125)       => (001.10001 | 1.53125)         
    1993 => 49,           -- (011111.001001 | 31.140625)    => (001.10001 | 1.53125)         
    1994 => 49,           -- (011111.001010 | 31.15625)     => (001.10001 | 1.53125)         
    1995 => 49,           -- (011111.001011 | 31.171875)    => (001.10001 | 1.53125)         
    1996 => 49,           -- (011111.001100 | 31.1875)      => (001.10001 | 1.53125)         
    1997 => 49,           -- (011111.001101 | 31.203125)    => (001.10001 | 1.53125)         
    1998 => 49,           -- (011111.001110 | 31.21875)     => (001.10001 | 1.53125)         
    1999 => 49,           -- (011111.001111 | 31.234375)    => (001.10001 | 1.53125)         
    2000 => 49,           -- (011111.010000 | 31.25)        => (001.10001 | 1.53125)         
    2001 => 49,           -- (011111.010001 | 31.265625)    => (001.10001 | 1.53125)         
    2002 => 49,           -- (011111.010010 | 31.28125)     => (001.10001 | 1.53125)         
    2003 => 49,           -- (011111.010011 | 31.296875)    => (001.10001 | 1.53125)         
    2004 => 49,           -- (011111.010100 | 31.3125)      => (001.10001 | 1.53125)         
    2005 => 49,           -- (011111.010101 | 31.328125)    => (001.10001 | 1.53125)         
    2006 => 49,           -- (011111.010110 | 31.34375)     => (001.10001 | 1.53125)         
    2007 => 49,           -- (011111.010111 | 31.359375)    => (001.10001 | 1.53125)         
    2008 => 49,           -- (011111.011000 | 31.375)       => (001.10001 | 1.53125)         
    2009 => 49,           -- (011111.011001 | 31.390625)    => (001.10001 | 1.53125)         
    2010 => 49,           -- (011111.011010 | 31.40625)     => (001.10001 | 1.53125)         
    2011 => 49,           -- (011111.011011 | 31.421875)    => (001.10001 | 1.53125)         
    2012 => 49,           -- (011111.011100 | 31.4375)      => (001.10001 | 1.53125)         
    2013 => 49,           -- (011111.011101 | 31.453125)    => (001.10001 | 1.53125)         
    2014 => 49,           -- (011111.011110 | 31.46875)     => (001.10001 | 1.53125)         
    2015 => 49,           -- (011111.011111 | 31.484375)    => (001.10001 | 1.53125)         
    2016 => 49,           -- (011111.100000 | 31.5)         => (001.10001 | 1.53125)         
    2017 => 49,           -- (011111.100001 | 31.515625)    => (001.10001 | 1.53125)         
    2018 => 49,           -- (011111.100010 | 31.53125)     => (001.10001 | 1.53125)         
    2019 => 49,           -- (011111.100011 | 31.546875)    => (001.10001 | 1.53125)         
    2020 => 49,           -- (011111.100100 | 31.5625)      => (001.10001 | 1.53125)         
    2021 => 49,           -- (011111.100101 | 31.578125)    => (001.10001 | 1.53125)         
    2022 => 49,           -- (011111.100110 | 31.59375)     => (001.10001 | 1.53125)         
    2023 => 49,           -- (011111.100111 | 31.609375)    => (001.10001 | 1.53125)         
    2024 => 49,           -- (011111.101000 | 31.625)       => (001.10001 | 1.53125)         
    2025 => 49,           -- (011111.101001 | 31.640625)    => (001.10001 | 1.53125)         
    2026 => 49,           -- (011111.101010 | 31.65625)     => (001.10001 | 1.53125)         
    2027 => 49,           -- (011111.101011 | 31.671875)    => (001.10001 | 1.53125)         
    2028 => 49,           -- (011111.101100 | 31.6875)      => (001.10001 | 1.53125)         
    2029 => 49,           -- (011111.101101 | 31.703125)    => (001.10001 | 1.53125)         
    2030 => 49,           -- (011111.101110 | 31.71875)     => (001.10001 | 1.53125)         
    2031 => 49,           -- (011111.101111 | 31.734375)    => (001.10001 | 1.53125)         
    2032 => 49,           -- (011111.110000 | 31.75)        => (001.10001 | 1.53125)         
    2033 => 49,           -- (011111.110001 | 31.765625)    => (001.10001 | 1.53125)         
    2034 => 49,           -- (011111.110010 | 31.78125)     => (001.10001 | 1.53125)         
    2035 => 49,           -- (011111.110011 | 31.796875)    => (001.10001 | 1.53125)         
    2036 => 49,           -- (011111.110100 | 31.8125)      => (001.10001 | 1.53125)         
    2037 => 49,           -- (011111.110101 | 31.828125)    => (001.10001 | 1.53125)         
    2038 => 49,           -- (011111.110110 | 31.84375)     => (001.10001 | 1.53125)         
    2039 => 49,           -- (011111.110111 | 31.859375)    => (001.10001 | 1.53125)         
    2040 => 49,           -- (011111.111000 | 31.875)       => (001.10001 | 1.53125)         
    2041 => 49,           -- (011111.111001 | 31.890625)    => (001.10001 | 1.53125)         
    2042 => 49,           -- (011111.111010 | 31.90625)     => (001.10001 | 1.53125)         
    2043 => 49,           -- (011111.111011 | 31.921875)    => (001.10001 | 1.53125)         
    2044 => 49,           -- (011111.111100 | 31.9375)      => (001.10001 | 1.53125)         
    2045 => 49,           -- (011111.111101 | 31.953125)    => (001.10001 | 1.53125)         
    2046 => 49,           -- (011111.111110 | 31.96875)     => (001.10001 | 1.53125)         
    2047 => 49,           -- (011111.111111 | 31.984375)    => (001.10001 | 1.53125)         
    2048 => 206,          -- (100000.000000 | -32.0)        => (110.01110 | -1.5625)         
    2049 => 206,          -- (100000.000001 | -31.984375)   => (110.01110 | -1.5625)         
    2050 => 206,          -- (100000.000010 | -31.96875)    => (110.01110 | -1.5625)         
    2051 => 206,          -- (100000.000011 | -31.953125)   => (110.01110 | -1.5625)         
    2052 => 206,          -- (100000.000100 | -31.9375)     => (110.01110 | -1.5625)         
    2053 => 206,          -- (100000.000101 | -31.921875)   => (110.01110 | -1.5625)         
    2054 => 206,          -- (100000.000110 | -31.90625)    => (110.01110 | -1.5625)         
    2055 => 206,          -- (100000.000111 | -31.890625)   => (110.01110 | -1.5625)         
    2056 => 206,          -- (100000.001000 | -31.875)      => (110.01110 | -1.5625)         
    2057 => 206,          -- (100000.001001 | -31.859375)   => (110.01110 | -1.5625)         
    2058 => 206,          -- (100000.001010 | -31.84375)    => (110.01110 | -1.5625)         
    2059 => 206,          -- (100000.001011 | -31.828125)   => (110.01110 | -1.5625)         
    2060 => 206,          -- (100000.001100 | -31.8125)     => (110.01110 | -1.5625)         
    2061 => 206,          -- (100000.001101 | -31.796875)   => (110.01110 | -1.5625)         
    2062 => 206,          -- (100000.001110 | -31.78125)    => (110.01110 | -1.5625)         
    2063 => 206,          -- (100000.001111 | -31.765625)   => (110.01110 | -1.5625)         
    2064 => 206,          -- (100000.010000 | -31.75)       => (110.01110 | -1.5625)         
    2065 => 206,          -- (100000.010001 | -31.734375)   => (110.01110 | -1.5625)         
    2066 => 206,          -- (100000.010010 | -31.71875)    => (110.01110 | -1.5625)         
    2067 => 206,          -- (100000.010011 | -31.703125)   => (110.01110 | -1.5625)         
    2068 => 206,          -- (100000.010100 | -31.6875)     => (110.01110 | -1.5625)         
    2069 => 206,          -- (100000.010101 | -31.671875)   => (110.01110 | -1.5625)         
    2070 => 206,          -- (100000.010110 | -31.65625)    => (110.01110 | -1.5625)         
    2071 => 206,          -- (100000.010111 | -31.640625)   => (110.01110 | -1.5625)         
    2072 => 206,          -- (100000.011000 | -31.625)      => (110.01110 | -1.5625)         
    2073 => 206,          -- (100000.011001 | -31.609375)   => (110.01110 | -1.5625)         
    2074 => 206,          -- (100000.011010 | -31.59375)    => (110.01110 | -1.5625)         
    2075 => 206,          -- (100000.011011 | -31.578125)   => (110.01110 | -1.5625)         
    2076 => 206,          -- (100000.011100 | -31.5625)     => (110.01110 | -1.5625)         
    2077 => 206,          -- (100000.011101 | -31.546875)   => (110.01110 | -1.5625)         
    2078 => 206,          -- (100000.011110 | -31.53125)    => (110.01110 | -1.5625)         
    2079 => 206,          -- (100000.011111 | -31.515625)   => (110.01110 | -1.5625)         
    2080 => 206,          -- (100000.100000 | -31.5)        => (110.01110 | -1.5625)         
    2081 => 206,          -- (100000.100001 | -31.484375)   => (110.01110 | -1.5625)         
    2082 => 206,          -- (100000.100010 | -31.46875)    => (110.01110 | -1.5625)         
    2083 => 206,          -- (100000.100011 | -31.453125)   => (110.01110 | -1.5625)         
    2084 => 206,          -- (100000.100100 | -31.4375)     => (110.01110 | -1.5625)         
    2085 => 206,          -- (100000.100101 | -31.421875)   => (110.01110 | -1.5625)         
    2086 => 206,          -- (100000.100110 | -31.40625)    => (110.01110 | -1.5625)         
    2087 => 206,          -- (100000.100111 | -31.390625)   => (110.01110 | -1.5625)         
    2088 => 206,          -- (100000.101000 | -31.375)      => (110.01110 | -1.5625)         
    2089 => 206,          -- (100000.101001 | -31.359375)   => (110.01110 | -1.5625)         
    2090 => 206,          -- (100000.101010 | -31.34375)    => (110.01110 | -1.5625)         
    2091 => 206,          -- (100000.101011 | -31.328125)   => (110.01110 | -1.5625)         
    2092 => 206,          -- (100000.101100 | -31.3125)     => (110.01110 | -1.5625)         
    2093 => 206,          -- (100000.101101 | -31.296875)   => (110.01110 | -1.5625)         
    2094 => 206,          -- (100000.101110 | -31.28125)    => (110.01110 | -1.5625)         
    2095 => 206,          -- (100000.101111 | -31.265625)   => (110.01110 | -1.5625)         
    2096 => 206,          -- (100000.110000 | -31.25)       => (110.01110 | -1.5625)         
    2097 => 206,          -- (100000.110001 | -31.234375)   => (110.01110 | -1.5625)         
    2098 => 206,          -- (100000.110010 | -31.21875)    => (110.01110 | -1.5625)         
    2099 => 206,          -- (100000.110011 | -31.203125)   => (110.01110 | -1.5625)         
    2100 => 206,          -- (100000.110100 | -31.1875)     => (110.01110 | -1.5625)         
    2101 => 206,          -- (100000.110101 | -31.171875)   => (110.01110 | -1.5625)         
    2102 => 206,          -- (100000.110110 | -31.15625)    => (110.01110 | -1.5625)         
    2103 => 206,          -- (100000.110111 | -31.140625)   => (110.01110 | -1.5625)         
    2104 => 206,          -- (100000.111000 | -31.125)      => (110.01110 | -1.5625)         
    2105 => 206,          -- (100000.111001 | -31.109375)   => (110.01110 | -1.5625)         
    2106 => 206,          -- (100000.111010 | -31.09375)    => (110.01110 | -1.5625)         
    2107 => 206,          -- (100000.111011 | -31.078125)   => (110.01110 | -1.5625)         
    2108 => 206,          -- (100000.111100 | -31.0625)     => (110.01110 | -1.5625)         
    2109 => 206,          -- (100000.111101 | -31.046875)   => (110.01110 | -1.5625)         
    2110 => 206,          -- (100000.111110 | -31.03125)    => (110.01110 | -1.5625)         
    2111 => 206,          -- (100000.111111 | -31.015625)   => (110.01110 | -1.5625)         
    2112 => 206,          -- (100001.000000 | -31.0)        => (110.01110 | -1.5625)         
    2113 => 206,          -- (100001.000001 | -30.984375)   => (110.01110 | -1.5625)         
    2114 => 206,          -- (100001.000010 | -30.96875)    => (110.01110 | -1.5625)         
    2115 => 206,          -- (100001.000011 | -30.953125)   => (110.01110 | -1.5625)         
    2116 => 206,          -- (100001.000100 | -30.9375)     => (110.01110 | -1.5625)         
    2117 => 206,          -- (100001.000101 | -30.921875)   => (110.01110 | -1.5625)         
    2118 => 206,          -- (100001.000110 | -30.90625)    => (110.01110 | -1.5625)         
    2119 => 206,          -- (100001.000111 | -30.890625)   => (110.01110 | -1.5625)         
    2120 => 206,          -- (100001.001000 | -30.875)      => (110.01110 | -1.5625)         
    2121 => 206,          -- (100001.001001 | -30.859375)   => (110.01110 | -1.5625)         
    2122 => 206,          -- (100001.001010 | -30.84375)    => (110.01110 | -1.5625)         
    2123 => 206,          -- (100001.001011 | -30.828125)   => (110.01110 | -1.5625)         
    2124 => 206,          -- (100001.001100 | -30.8125)     => (110.01110 | -1.5625)         
    2125 => 206,          -- (100001.001101 | -30.796875)   => (110.01110 | -1.5625)         
    2126 => 206,          -- (100001.001110 | -30.78125)    => (110.01110 | -1.5625)         
    2127 => 206,          -- (100001.001111 | -30.765625)   => (110.01110 | -1.5625)         
    2128 => 206,          -- (100001.010000 | -30.75)       => (110.01110 | -1.5625)         
    2129 => 206,          -- (100001.010001 | -30.734375)   => (110.01110 | -1.5625)         
    2130 => 206,          -- (100001.010010 | -30.71875)    => (110.01110 | -1.5625)         
    2131 => 206,          -- (100001.010011 | -30.703125)   => (110.01110 | -1.5625)         
    2132 => 206,          -- (100001.010100 | -30.6875)     => (110.01110 | -1.5625)         
    2133 => 206,          -- (100001.010101 | -30.671875)   => (110.01110 | -1.5625)         
    2134 => 206,          -- (100001.010110 | -30.65625)    => (110.01110 | -1.5625)         
    2135 => 206,          -- (100001.010111 | -30.640625)   => (110.01110 | -1.5625)         
    2136 => 206,          -- (100001.011000 | -30.625)      => (110.01110 | -1.5625)         
    2137 => 206,          -- (100001.011001 | -30.609375)   => (110.01110 | -1.5625)         
    2138 => 206,          -- (100001.011010 | -30.59375)    => (110.01110 | -1.5625)         
    2139 => 206,          -- (100001.011011 | -30.578125)   => (110.01110 | -1.5625)         
    2140 => 206,          -- (100001.011100 | -30.5625)     => (110.01110 | -1.5625)         
    2141 => 206,          -- (100001.011101 | -30.546875)   => (110.01110 | -1.5625)         
    2142 => 206,          -- (100001.011110 | -30.53125)    => (110.01110 | -1.5625)         
    2143 => 206,          -- (100001.011111 | -30.515625)   => (110.01110 | -1.5625)         
    2144 => 206,          -- (100001.100000 | -30.5)        => (110.01110 | -1.5625)         
    2145 => 206,          -- (100001.100001 | -30.484375)   => (110.01110 | -1.5625)         
    2146 => 206,          -- (100001.100010 | -30.46875)    => (110.01110 | -1.5625)         
    2147 => 206,          -- (100001.100011 | -30.453125)   => (110.01110 | -1.5625)         
    2148 => 206,          -- (100001.100100 | -30.4375)     => (110.01110 | -1.5625)         
    2149 => 206,          -- (100001.100101 | -30.421875)   => (110.01110 | -1.5625)         
    2150 => 206,          -- (100001.100110 | -30.40625)    => (110.01110 | -1.5625)         
    2151 => 206,          -- (100001.100111 | -30.390625)   => (110.01110 | -1.5625)         
    2152 => 206,          -- (100001.101000 | -30.375)      => (110.01110 | -1.5625)         
    2153 => 206,          -- (100001.101001 | -30.359375)   => (110.01110 | -1.5625)         
    2154 => 206,          -- (100001.101010 | -30.34375)    => (110.01110 | -1.5625)         
    2155 => 206,          -- (100001.101011 | -30.328125)   => (110.01110 | -1.5625)         
    2156 => 206,          -- (100001.101100 | -30.3125)     => (110.01110 | -1.5625)         
    2157 => 206,          -- (100001.101101 | -30.296875)   => (110.01110 | -1.5625)         
    2158 => 206,          -- (100001.101110 | -30.28125)    => (110.01110 | -1.5625)         
    2159 => 206,          -- (100001.101111 | -30.265625)   => (110.01110 | -1.5625)         
    2160 => 206,          -- (100001.110000 | -30.25)       => (110.01110 | -1.5625)         
    2161 => 206,          -- (100001.110001 | -30.234375)   => (110.01110 | -1.5625)         
    2162 => 206,          -- (100001.110010 | -30.21875)    => (110.01110 | -1.5625)         
    2163 => 206,          -- (100001.110011 | -30.203125)   => (110.01110 | -1.5625)         
    2164 => 206,          -- (100001.110100 | -30.1875)     => (110.01110 | -1.5625)         
    2165 => 206,          -- (100001.110101 | -30.171875)   => (110.01110 | -1.5625)         
    2166 => 206,          -- (100001.110110 | -30.15625)    => (110.01110 | -1.5625)         
    2167 => 206,          -- (100001.110111 | -30.140625)   => (110.01110 | -1.5625)         
    2168 => 206,          -- (100001.111000 | -30.125)      => (110.01110 | -1.5625)         
    2169 => 206,          -- (100001.111001 | -30.109375)   => (110.01110 | -1.5625)         
    2170 => 206,          -- (100001.111010 | -30.09375)    => (110.01110 | -1.5625)         
    2171 => 206,          -- (100001.111011 | -30.078125)   => (110.01110 | -1.5625)         
    2172 => 206,          -- (100001.111100 | -30.0625)     => (110.01110 | -1.5625)         
    2173 => 206,          -- (100001.111101 | -30.046875)   => (110.01110 | -1.5625)         
    2174 => 206,          -- (100001.111110 | -30.03125)    => (110.01110 | -1.5625)         
    2175 => 206,          -- (100001.111111 | -30.015625)   => (110.01110 | -1.5625)         
    2176 => 206,          -- (100010.000000 | -30.0)        => (110.01110 | -1.5625)         
    2177 => 206,          -- (100010.000001 | -29.984375)   => (110.01110 | -1.5625)         
    2178 => 206,          -- (100010.000010 | -29.96875)    => (110.01110 | -1.5625)         
    2179 => 206,          -- (100010.000011 | -29.953125)   => (110.01110 | -1.5625)         
    2180 => 206,          -- (100010.000100 | -29.9375)     => (110.01110 | -1.5625)         
    2181 => 206,          -- (100010.000101 | -29.921875)   => (110.01110 | -1.5625)         
    2182 => 206,          -- (100010.000110 | -29.90625)    => (110.01110 | -1.5625)         
    2183 => 206,          -- (100010.000111 | -29.890625)   => (110.01110 | -1.5625)         
    2184 => 206,          -- (100010.001000 | -29.875)      => (110.01110 | -1.5625)         
    2185 => 206,          -- (100010.001001 | -29.859375)   => (110.01110 | -1.5625)         
    2186 => 206,          -- (100010.001010 | -29.84375)    => (110.01110 | -1.5625)         
    2187 => 206,          -- (100010.001011 | -29.828125)   => (110.01110 | -1.5625)         
    2188 => 206,          -- (100010.001100 | -29.8125)     => (110.01110 | -1.5625)         
    2189 => 206,          -- (100010.001101 | -29.796875)   => (110.01110 | -1.5625)         
    2190 => 206,          -- (100010.001110 | -29.78125)    => (110.01110 | -1.5625)         
    2191 => 206,          -- (100010.001111 | -29.765625)   => (110.01110 | -1.5625)         
    2192 => 206,          -- (100010.010000 | -29.75)       => (110.01110 | -1.5625)         
    2193 => 206,          -- (100010.010001 | -29.734375)   => (110.01110 | -1.5625)         
    2194 => 206,          -- (100010.010010 | -29.71875)    => (110.01110 | -1.5625)         
    2195 => 206,          -- (100010.010011 | -29.703125)   => (110.01110 | -1.5625)         
    2196 => 206,          -- (100010.010100 | -29.6875)     => (110.01110 | -1.5625)         
    2197 => 206,          -- (100010.010101 | -29.671875)   => (110.01110 | -1.5625)         
    2198 => 206,          -- (100010.010110 | -29.65625)    => (110.01110 | -1.5625)         
    2199 => 206,          -- (100010.010111 | -29.640625)   => (110.01110 | -1.5625)         
    2200 => 206,          -- (100010.011000 | -29.625)      => (110.01110 | -1.5625)         
    2201 => 206,          -- (100010.011001 | -29.609375)   => (110.01110 | -1.5625)         
    2202 => 206,          -- (100010.011010 | -29.59375)    => (110.01110 | -1.5625)         
    2203 => 206,          -- (100010.011011 | -29.578125)   => (110.01110 | -1.5625)         
    2204 => 206,          -- (100010.011100 | -29.5625)     => (110.01110 | -1.5625)         
    2205 => 206,          -- (100010.011101 | -29.546875)   => (110.01110 | -1.5625)         
    2206 => 206,          -- (100010.011110 | -29.53125)    => (110.01110 | -1.5625)         
    2207 => 206,          -- (100010.011111 | -29.515625)   => (110.01110 | -1.5625)         
    2208 => 206,          -- (100010.100000 | -29.5)        => (110.01110 | -1.5625)         
    2209 => 206,          -- (100010.100001 | -29.484375)   => (110.01110 | -1.5625)         
    2210 => 206,          -- (100010.100010 | -29.46875)    => (110.01110 | -1.5625)         
    2211 => 206,          -- (100010.100011 | -29.453125)   => (110.01110 | -1.5625)         
    2212 => 206,          -- (100010.100100 | -29.4375)     => (110.01110 | -1.5625)         
    2213 => 206,          -- (100010.100101 | -29.421875)   => (110.01110 | -1.5625)         
    2214 => 206,          -- (100010.100110 | -29.40625)    => (110.01110 | -1.5625)         
    2215 => 206,          -- (100010.100111 | -29.390625)   => (110.01110 | -1.5625)         
    2216 => 206,          -- (100010.101000 | -29.375)      => (110.01110 | -1.5625)         
    2217 => 206,          -- (100010.101001 | -29.359375)   => (110.01110 | -1.5625)         
    2218 => 206,          -- (100010.101010 | -29.34375)    => (110.01110 | -1.5625)         
    2219 => 206,          -- (100010.101011 | -29.328125)   => (110.01110 | -1.5625)         
    2220 => 206,          -- (100010.101100 | -29.3125)     => (110.01110 | -1.5625)         
    2221 => 206,          -- (100010.101101 | -29.296875)   => (110.01110 | -1.5625)         
    2222 => 206,          -- (100010.101110 | -29.28125)    => (110.01110 | -1.5625)         
    2223 => 206,          -- (100010.101111 | -29.265625)   => (110.01110 | -1.5625)         
    2224 => 206,          -- (100010.110000 | -29.25)       => (110.01110 | -1.5625)         
    2225 => 206,          -- (100010.110001 | -29.234375)   => (110.01110 | -1.5625)         
    2226 => 206,          -- (100010.110010 | -29.21875)    => (110.01110 | -1.5625)         
    2227 => 206,          -- (100010.110011 | -29.203125)   => (110.01110 | -1.5625)         
    2228 => 206,          -- (100010.110100 | -29.1875)     => (110.01110 | -1.5625)         
    2229 => 206,          -- (100010.110101 | -29.171875)   => (110.01110 | -1.5625)         
    2230 => 206,          -- (100010.110110 | -29.15625)    => (110.01110 | -1.5625)         
    2231 => 206,          -- (100010.110111 | -29.140625)   => (110.01110 | -1.5625)         
    2232 => 206,          -- (100010.111000 | -29.125)      => (110.01110 | -1.5625)         
    2233 => 206,          -- (100010.111001 | -29.109375)   => (110.01110 | -1.5625)         
    2234 => 206,          -- (100010.111010 | -29.09375)    => (110.01110 | -1.5625)         
    2235 => 206,          -- (100010.111011 | -29.078125)   => (110.01110 | -1.5625)         
    2236 => 206,          -- (100010.111100 | -29.0625)     => (110.01110 | -1.5625)         
    2237 => 206,          -- (100010.111101 | -29.046875)   => (110.01110 | -1.5625)         
    2238 => 206,          -- (100010.111110 | -29.03125)    => (110.01110 | -1.5625)         
    2239 => 206,          -- (100010.111111 | -29.015625)   => (110.01110 | -1.5625)         
    2240 => 206,          -- (100011.000000 | -29.0)        => (110.01110 | -1.5625)         
    2241 => 206,          -- (100011.000001 | -28.984375)   => (110.01110 | -1.5625)         
    2242 => 206,          -- (100011.000010 | -28.96875)    => (110.01110 | -1.5625)         
    2243 => 206,          -- (100011.000011 | -28.953125)   => (110.01110 | -1.5625)         
    2244 => 206,          -- (100011.000100 | -28.9375)     => (110.01110 | -1.5625)         
    2245 => 206,          -- (100011.000101 | -28.921875)   => (110.01110 | -1.5625)         
    2246 => 206,          -- (100011.000110 | -28.90625)    => (110.01110 | -1.5625)         
    2247 => 206,          -- (100011.000111 | -28.890625)   => (110.01110 | -1.5625)         
    2248 => 206,          -- (100011.001000 | -28.875)      => (110.01110 | -1.5625)         
    2249 => 206,          -- (100011.001001 | -28.859375)   => (110.01110 | -1.5625)         
    2250 => 206,          -- (100011.001010 | -28.84375)    => (110.01110 | -1.5625)         
    2251 => 206,          -- (100011.001011 | -28.828125)   => (110.01110 | -1.5625)         
    2252 => 206,          -- (100011.001100 | -28.8125)     => (110.01110 | -1.5625)         
    2253 => 206,          -- (100011.001101 | -28.796875)   => (110.01110 | -1.5625)         
    2254 => 206,          -- (100011.001110 | -28.78125)    => (110.01110 | -1.5625)         
    2255 => 206,          -- (100011.001111 | -28.765625)   => (110.01110 | -1.5625)         
    2256 => 206,          -- (100011.010000 | -28.75)       => (110.01110 | -1.5625)         
    2257 => 206,          -- (100011.010001 | -28.734375)   => (110.01110 | -1.5625)         
    2258 => 206,          -- (100011.010010 | -28.71875)    => (110.01110 | -1.5625)         
    2259 => 206,          -- (100011.010011 | -28.703125)   => (110.01110 | -1.5625)         
    2260 => 206,          -- (100011.010100 | -28.6875)     => (110.01110 | -1.5625)         
    2261 => 206,          -- (100011.010101 | -28.671875)   => (110.01110 | -1.5625)         
    2262 => 206,          -- (100011.010110 | -28.65625)    => (110.01110 | -1.5625)         
    2263 => 206,          -- (100011.010111 | -28.640625)   => (110.01110 | -1.5625)         
    2264 => 206,          -- (100011.011000 | -28.625)      => (110.01110 | -1.5625)         
    2265 => 206,          -- (100011.011001 | -28.609375)   => (110.01110 | -1.5625)         
    2266 => 206,          -- (100011.011010 | -28.59375)    => (110.01110 | -1.5625)         
    2267 => 206,          -- (100011.011011 | -28.578125)   => (110.01110 | -1.5625)         
    2268 => 206,          -- (100011.011100 | -28.5625)     => (110.01110 | -1.5625)         
    2269 => 206,          -- (100011.011101 | -28.546875)   => (110.01110 | -1.5625)         
    2270 => 206,          -- (100011.011110 | -28.53125)    => (110.01110 | -1.5625)         
    2271 => 206,          -- (100011.011111 | -28.515625)   => (110.01110 | -1.5625)         
    2272 => 206,          -- (100011.100000 | -28.5)        => (110.01110 | -1.5625)         
    2273 => 206,          -- (100011.100001 | -28.484375)   => (110.01110 | -1.5625)         
    2274 => 206,          -- (100011.100010 | -28.46875)    => (110.01110 | -1.5625)         
    2275 => 206,          -- (100011.100011 | -28.453125)   => (110.01110 | -1.5625)         
    2276 => 206,          -- (100011.100100 | -28.4375)     => (110.01110 | -1.5625)         
    2277 => 206,          -- (100011.100101 | -28.421875)   => (110.01110 | -1.5625)         
    2278 => 206,          -- (100011.100110 | -28.40625)    => (110.01110 | -1.5625)         
    2279 => 206,          -- (100011.100111 | -28.390625)   => (110.01110 | -1.5625)         
    2280 => 206,          -- (100011.101000 | -28.375)      => (110.01110 | -1.5625)         
    2281 => 206,          -- (100011.101001 | -28.359375)   => (110.01110 | -1.5625)         
    2282 => 206,          -- (100011.101010 | -28.34375)    => (110.01110 | -1.5625)         
    2283 => 206,          -- (100011.101011 | -28.328125)   => (110.01110 | -1.5625)         
    2284 => 206,          -- (100011.101100 | -28.3125)     => (110.01110 | -1.5625)         
    2285 => 206,          -- (100011.101101 | -28.296875)   => (110.01110 | -1.5625)         
    2286 => 206,          -- (100011.101110 | -28.28125)    => (110.01110 | -1.5625)         
    2287 => 206,          -- (100011.101111 | -28.265625)   => (110.01110 | -1.5625)         
    2288 => 206,          -- (100011.110000 | -28.25)       => (110.01110 | -1.5625)         
    2289 => 206,          -- (100011.110001 | -28.234375)   => (110.01110 | -1.5625)         
    2290 => 206,          -- (100011.110010 | -28.21875)    => (110.01110 | -1.5625)         
    2291 => 206,          -- (100011.110011 | -28.203125)   => (110.01110 | -1.5625)         
    2292 => 206,          -- (100011.110100 | -28.1875)     => (110.01110 | -1.5625)         
    2293 => 206,          -- (100011.110101 | -28.171875)   => (110.01110 | -1.5625)         
    2294 => 206,          -- (100011.110110 | -28.15625)    => (110.01110 | -1.5625)         
    2295 => 206,          -- (100011.110111 | -28.140625)   => (110.01110 | -1.5625)         
    2296 => 206,          -- (100011.111000 | -28.125)      => (110.01110 | -1.5625)         
    2297 => 206,          -- (100011.111001 | -28.109375)   => (110.01110 | -1.5625)         
    2298 => 206,          -- (100011.111010 | -28.09375)    => (110.01110 | -1.5625)         
    2299 => 206,          -- (100011.111011 | -28.078125)   => (110.01110 | -1.5625)         
    2300 => 206,          -- (100011.111100 | -28.0625)     => (110.01110 | -1.5625)         
    2301 => 206,          -- (100011.111101 | -28.046875)   => (110.01110 | -1.5625)         
    2302 => 206,          -- (100011.111110 | -28.03125)    => (110.01110 | -1.5625)         
    2303 => 206,          -- (100011.111111 | -28.015625)   => (110.01110 | -1.5625)         
    2304 => 206,          -- (100100.000000 | -28.0)        => (110.01110 | -1.5625)         
    2305 => 206,          -- (100100.000001 | -27.984375)   => (110.01110 | -1.5625)         
    2306 => 206,          -- (100100.000010 | -27.96875)    => (110.01110 | -1.5625)         
    2307 => 206,          -- (100100.000011 | -27.953125)   => (110.01110 | -1.5625)         
    2308 => 206,          -- (100100.000100 | -27.9375)     => (110.01110 | -1.5625)         
    2309 => 206,          -- (100100.000101 | -27.921875)   => (110.01110 | -1.5625)         
    2310 => 206,          -- (100100.000110 | -27.90625)    => (110.01110 | -1.5625)         
    2311 => 206,          -- (100100.000111 | -27.890625)   => (110.01110 | -1.5625)         
    2312 => 206,          -- (100100.001000 | -27.875)      => (110.01110 | -1.5625)         
    2313 => 206,          -- (100100.001001 | -27.859375)   => (110.01110 | -1.5625)         
    2314 => 206,          -- (100100.001010 | -27.84375)    => (110.01110 | -1.5625)         
    2315 => 206,          -- (100100.001011 | -27.828125)   => (110.01110 | -1.5625)         
    2316 => 206,          -- (100100.001100 | -27.8125)     => (110.01110 | -1.5625)         
    2317 => 206,          -- (100100.001101 | -27.796875)   => (110.01110 | -1.5625)         
    2318 => 206,          -- (100100.001110 | -27.78125)    => (110.01110 | -1.5625)         
    2319 => 206,          -- (100100.001111 | -27.765625)   => (110.01110 | -1.5625)         
    2320 => 206,          -- (100100.010000 | -27.75)       => (110.01110 | -1.5625)         
    2321 => 206,          -- (100100.010001 | -27.734375)   => (110.01110 | -1.5625)         
    2322 => 206,          -- (100100.010010 | -27.71875)    => (110.01110 | -1.5625)         
    2323 => 206,          -- (100100.010011 | -27.703125)   => (110.01110 | -1.5625)         
    2324 => 206,          -- (100100.010100 | -27.6875)     => (110.01110 | -1.5625)         
    2325 => 206,          -- (100100.010101 | -27.671875)   => (110.01110 | -1.5625)         
    2326 => 206,          -- (100100.010110 | -27.65625)    => (110.01110 | -1.5625)         
    2327 => 206,          -- (100100.010111 | -27.640625)   => (110.01110 | -1.5625)         
    2328 => 206,          -- (100100.011000 | -27.625)      => (110.01110 | -1.5625)         
    2329 => 206,          -- (100100.011001 | -27.609375)   => (110.01110 | -1.5625)         
    2330 => 206,          -- (100100.011010 | -27.59375)    => (110.01110 | -1.5625)         
    2331 => 206,          -- (100100.011011 | -27.578125)   => (110.01110 | -1.5625)         
    2332 => 206,          -- (100100.011100 | -27.5625)     => (110.01110 | -1.5625)         
    2333 => 206,          -- (100100.011101 | -27.546875)   => (110.01110 | -1.5625)         
    2334 => 206,          -- (100100.011110 | -27.53125)    => (110.01110 | -1.5625)         
    2335 => 206,          -- (100100.011111 | -27.515625)   => (110.01110 | -1.5625)         
    2336 => 206,          -- (100100.100000 | -27.5)        => (110.01110 | -1.5625)         
    2337 => 206,          -- (100100.100001 | -27.484375)   => (110.01110 | -1.5625)         
    2338 => 206,          -- (100100.100010 | -27.46875)    => (110.01110 | -1.5625)         
    2339 => 206,          -- (100100.100011 | -27.453125)   => (110.01110 | -1.5625)         
    2340 => 206,          -- (100100.100100 | -27.4375)     => (110.01110 | -1.5625)         
    2341 => 206,          -- (100100.100101 | -27.421875)   => (110.01110 | -1.5625)         
    2342 => 206,          -- (100100.100110 | -27.40625)    => (110.01110 | -1.5625)         
    2343 => 206,          -- (100100.100111 | -27.390625)   => (110.01110 | -1.5625)         
    2344 => 206,          -- (100100.101000 | -27.375)      => (110.01110 | -1.5625)         
    2345 => 206,          -- (100100.101001 | -27.359375)   => (110.01110 | -1.5625)         
    2346 => 206,          -- (100100.101010 | -27.34375)    => (110.01110 | -1.5625)         
    2347 => 206,          -- (100100.101011 | -27.328125)   => (110.01110 | -1.5625)         
    2348 => 206,          -- (100100.101100 | -27.3125)     => (110.01110 | -1.5625)         
    2349 => 206,          -- (100100.101101 | -27.296875)   => (110.01110 | -1.5625)         
    2350 => 206,          -- (100100.101110 | -27.28125)    => (110.01110 | -1.5625)         
    2351 => 206,          -- (100100.101111 | -27.265625)   => (110.01110 | -1.5625)         
    2352 => 206,          -- (100100.110000 | -27.25)       => (110.01110 | -1.5625)         
    2353 => 206,          -- (100100.110001 | -27.234375)   => (110.01110 | -1.5625)         
    2354 => 206,          -- (100100.110010 | -27.21875)    => (110.01110 | -1.5625)         
    2355 => 206,          -- (100100.110011 | -27.203125)   => (110.01110 | -1.5625)         
    2356 => 206,          -- (100100.110100 | -27.1875)     => (110.01110 | -1.5625)         
    2357 => 206,          -- (100100.110101 | -27.171875)   => (110.01110 | -1.5625)         
    2358 => 206,          -- (100100.110110 | -27.15625)    => (110.01110 | -1.5625)         
    2359 => 206,          -- (100100.110111 | -27.140625)   => (110.01110 | -1.5625)         
    2360 => 206,          -- (100100.111000 | -27.125)      => (110.01110 | -1.5625)         
    2361 => 206,          -- (100100.111001 | -27.109375)   => (110.01110 | -1.5625)         
    2362 => 206,          -- (100100.111010 | -27.09375)    => (110.01110 | -1.5625)         
    2363 => 206,          -- (100100.111011 | -27.078125)   => (110.01110 | -1.5625)         
    2364 => 206,          -- (100100.111100 | -27.0625)     => (110.01110 | -1.5625)         
    2365 => 206,          -- (100100.111101 | -27.046875)   => (110.01110 | -1.5625)         
    2366 => 206,          -- (100100.111110 | -27.03125)    => (110.01110 | -1.5625)         
    2367 => 206,          -- (100100.111111 | -27.015625)   => (110.01110 | -1.5625)         
    2368 => 206,          -- (100101.000000 | -27.0)        => (110.01110 | -1.5625)         
    2369 => 206,          -- (100101.000001 | -26.984375)   => (110.01110 | -1.5625)         
    2370 => 206,          -- (100101.000010 | -26.96875)    => (110.01110 | -1.5625)         
    2371 => 206,          -- (100101.000011 | -26.953125)   => (110.01110 | -1.5625)         
    2372 => 206,          -- (100101.000100 | -26.9375)     => (110.01110 | -1.5625)         
    2373 => 206,          -- (100101.000101 | -26.921875)   => (110.01110 | -1.5625)         
    2374 => 206,          -- (100101.000110 | -26.90625)    => (110.01110 | -1.5625)         
    2375 => 206,          -- (100101.000111 | -26.890625)   => (110.01110 | -1.5625)         
    2376 => 206,          -- (100101.001000 | -26.875)      => (110.01110 | -1.5625)         
    2377 => 206,          -- (100101.001001 | -26.859375)   => (110.01110 | -1.5625)         
    2378 => 206,          -- (100101.001010 | -26.84375)    => (110.01110 | -1.5625)         
    2379 => 206,          -- (100101.001011 | -26.828125)   => (110.01110 | -1.5625)         
    2380 => 206,          -- (100101.001100 | -26.8125)     => (110.01110 | -1.5625)         
    2381 => 206,          -- (100101.001101 | -26.796875)   => (110.01110 | -1.5625)         
    2382 => 206,          -- (100101.001110 | -26.78125)    => (110.01110 | -1.5625)         
    2383 => 206,          -- (100101.001111 | -26.765625)   => (110.01110 | -1.5625)         
    2384 => 206,          -- (100101.010000 | -26.75)       => (110.01110 | -1.5625)         
    2385 => 206,          -- (100101.010001 | -26.734375)   => (110.01110 | -1.5625)         
    2386 => 206,          -- (100101.010010 | -26.71875)    => (110.01110 | -1.5625)         
    2387 => 206,          -- (100101.010011 | -26.703125)   => (110.01110 | -1.5625)         
    2388 => 206,          -- (100101.010100 | -26.6875)     => (110.01110 | -1.5625)         
    2389 => 206,          -- (100101.010101 | -26.671875)   => (110.01110 | -1.5625)         
    2390 => 206,          -- (100101.010110 | -26.65625)    => (110.01110 | -1.5625)         
    2391 => 206,          -- (100101.010111 | -26.640625)   => (110.01110 | -1.5625)         
    2392 => 206,          -- (100101.011000 | -26.625)      => (110.01110 | -1.5625)         
    2393 => 206,          -- (100101.011001 | -26.609375)   => (110.01110 | -1.5625)         
    2394 => 206,          -- (100101.011010 | -26.59375)    => (110.01110 | -1.5625)         
    2395 => 206,          -- (100101.011011 | -26.578125)   => (110.01110 | -1.5625)         
    2396 => 206,          -- (100101.011100 | -26.5625)     => (110.01110 | -1.5625)         
    2397 => 206,          -- (100101.011101 | -26.546875)   => (110.01110 | -1.5625)         
    2398 => 206,          -- (100101.011110 | -26.53125)    => (110.01110 | -1.5625)         
    2399 => 206,          -- (100101.011111 | -26.515625)   => (110.01110 | -1.5625)         
    2400 => 206,          -- (100101.100000 | -26.5)        => (110.01110 | -1.5625)         
    2401 => 206,          -- (100101.100001 | -26.484375)   => (110.01110 | -1.5625)         
    2402 => 206,          -- (100101.100010 | -26.46875)    => (110.01110 | -1.5625)         
    2403 => 206,          -- (100101.100011 | -26.453125)   => (110.01110 | -1.5625)         
    2404 => 206,          -- (100101.100100 | -26.4375)     => (110.01110 | -1.5625)         
    2405 => 206,          -- (100101.100101 | -26.421875)   => (110.01110 | -1.5625)         
    2406 => 206,          -- (100101.100110 | -26.40625)    => (110.01110 | -1.5625)         
    2407 => 206,          -- (100101.100111 | -26.390625)   => (110.01110 | -1.5625)         
    2408 => 206,          -- (100101.101000 | -26.375)      => (110.01110 | -1.5625)         
    2409 => 206,          -- (100101.101001 | -26.359375)   => (110.01110 | -1.5625)         
    2410 => 206,          -- (100101.101010 | -26.34375)    => (110.01110 | -1.5625)         
    2411 => 206,          -- (100101.101011 | -26.328125)   => (110.01110 | -1.5625)         
    2412 => 206,          -- (100101.101100 | -26.3125)     => (110.01110 | -1.5625)         
    2413 => 206,          -- (100101.101101 | -26.296875)   => (110.01110 | -1.5625)         
    2414 => 206,          -- (100101.101110 | -26.28125)    => (110.01110 | -1.5625)         
    2415 => 206,          -- (100101.101111 | -26.265625)   => (110.01110 | -1.5625)         
    2416 => 206,          -- (100101.110000 | -26.25)       => (110.01110 | -1.5625)         
    2417 => 206,          -- (100101.110001 | -26.234375)   => (110.01110 | -1.5625)         
    2418 => 206,          -- (100101.110010 | -26.21875)    => (110.01110 | -1.5625)         
    2419 => 206,          -- (100101.110011 | -26.203125)   => (110.01110 | -1.5625)         
    2420 => 206,          -- (100101.110100 | -26.1875)     => (110.01110 | -1.5625)         
    2421 => 206,          -- (100101.110101 | -26.171875)   => (110.01110 | -1.5625)         
    2422 => 206,          -- (100101.110110 | -26.15625)    => (110.01110 | -1.5625)         
    2423 => 206,          -- (100101.110111 | -26.140625)   => (110.01110 | -1.5625)         
    2424 => 206,          -- (100101.111000 | -26.125)      => (110.01110 | -1.5625)         
    2425 => 206,          -- (100101.111001 | -26.109375)   => (110.01110 | -1.5625)         
    2426 => 206,          -- (100101.111010 | -26.09375)    => (110.01110 | -1.5625)         
    2427 => 206,          -- (100101.111011 | -26.078125)   => (110.01110 | -1.5625)         
    2428 => 206,          -- (100101.111100 | -26.0625)     => (110.01110 | -1.5625)         
    2429 => 206,          -- (100101.111101 | -26.046875)   => (110.01110 | -1.5625)         
    2430 => 206,          -- (100101.111110 | -26.03125)    => (110.01110 | -1.5625)         
    2431 => 206,          -- (100101.111111 | -26.015625)   => (110.01110 | -1.5625)         
    2432 => 206,          -- (100110.000000 | -26.0)        => (110.01110 | -1.5625)         
    2433 => 206,          -- (100110.000001 | -25.984375)   => (110.01110 | -1.5625)         
    2434 => 206,          -- (100110.000010 | -25.96875)    => (110.01110 | -1.5625)         
    2435 => 206,          -- (100110.000011 | -25.953125)   => (110.01110 | -1.5625)         
    2436 => 206,          -- (100110.000100 | -25.9375)     => (110.01110 | -1.5625)         
    2437 => 206,          -- (100110.000101 | -25.921875)   => (110.01110 | -1.5625)         
    2438 => 206,          -- (100110.000110 | -25.90625)    => (110.01110 | -1.5625)         
    2439 => 206,          -- (100110.000111 | -25.890625)   => (110.01110 | -1.5625)         
    2440 => 206,          -- (100110.001000 | -25.875)      => (110.01110 | -1.5625)         
    2441 => 206,          -- (100110.001001 | -25.859375)   => (110.01110 | -1.5625)         
    2442 => 206,          -- (100110.001010 | -25.84375)    => (110.01110 | -1.5625)         
    2443 => 206,          -- (100110.001011 | -25.828125)   => (110.01110 | -1.5625)         
    2444 => 206,          -- (100110.001100 | -25.8125)     => (110.01110 | -1.5625)         
    2445 => 206,          -- (100110.001101 | -25.796875)   => (110.01110 | -1.5625)         
    2446 => 206,          -- (100110.001110 | -25.78125)    => (110.01110 | -1.5625)         
    2447 => 206,          -- (100110.001111 | -25.765625)   => (110.01110 | -1.5625)         
    2448 => 206,          -- (100110.010000 | -25.75)       => (110.01110 | -1.5625)         
    2449 => 206,          -- (100110.010001 | -25.734375)   => (110.01110 | -1.5625)         
    2450 => 206,          -- (100110.010010 | -25.71875)    => (110.01110 | -1.5625)         
    2451 => 206,          -- (100110.010011 | -25.703125)   => (110.01110 | -1.5625)         
    2452 => 206,          -- (100110.010100 | -25.6875)     => (110.01110 | -1.5625)         
    2453 => 206,          -- (100110.010101 | -25.671875)   => (110.01110 | -1.5625)         
    2454 => 206,          -- (100110.010110 | -25.65625)    => (110.01110 | -1.5625)         
    2455 => 206,          -- (100110.010111 | -25.640625)   => (110.01110 | -1.5625)         
    2456 => 206,          -- (100110.011000 | -25.625)      => (110.01110 | -1.5625)         
    2457 => 206,          -- (100110.011001 | -25.609375)   => (110.01110 | -1.5625)         
    2458 => 206,          -- (100110.011010 | -25.59375)    => (110.01110 | -1.5625)         
    2459 => 206,          -- (100110.011011 | -25.578125)   => (110.01110 | -1.5625)         
    2460 => 206,          -- (100110.011100 | -25.5625)     => (110.01110 | -1.5625)         
    2461 => 206,          -- (100110.011101 | -25.546875)   => (110.01110 | -1.5625)         
    2462 => 206,          -- (100110.011110 | -25.53125)    => (110.01110 | -1.5625)         
    2463 => 206,          -- (100110.011111 | -25.515625)   => (110.01110 | -1.5625)         
    2464 => 206,          -- (100110.100000 | -25.5)        => (110.01110 | -1.5625)         
    2465 => 206,          -- (100110.100001 | -25.484375)   => (110.01110 | -1.5625)         
    2466 => 206,          -- (100110.100010 | -25.46875)    => (110.01110 | -1.5625)         
    2467 => 206,          -- (100110.100011 | -25.453125)   => (110.01110 | -1.5625)         
    2468 => 206,          -- (100110.100100 | -25.4375)     => (110.01110 | -1.5625)         
    2469 => 206,          -- (100110.100101 | -25.421875)   => (110.01110 | -1.5625)         
    2470 => 206,          -- (100110.100110 | -25.40625)    => (110.01110 | -1.5625)         
    2471 => 206,          -- (100110.100111 | -25.390625)   => (110.01110 | -1.5625)         
    2472 => 206,          -- (100110.101000 | -25.375)      => (110.01110 | -1.5625)         
    2473 => 206,          -- (100110.101001 | -25.359375)   => (110.01110 | -1.5625)         
    2474 => 206,          -- (100110.101010 | -25.34375)    => (110.01110 | -1.5625)         
    2475 => 206,          -- (100110.101011 | -25.328125)   => (110.01110 | -1.5625)         
    2476 => 206,          -- (100110.101100 | -25.3125)     => (110.01110 | -1.5625)         
    2477 => 206,          -- (100110.101101 | -25.296875)   => (110.01110 | -1.5625)         
    2478 => 206,          -- (100110.101110 | -25.28125)    => (110.01110 | -1.5625)         
    2479 => 207,          -- (100110.101111 | -25.265625)   => (110.01111 | -1.53125)        
    2480 => 207,          -- (100110.110000 | -25.25)       => (110.01111 | -1.53125)        
    2481 => 207,          -- (100110.110001 | -25.234375)   => (110.01111 | -1.53125)        
    2482 => 207,          -- (100110.110010 | -25.21875)    => (110.01111 | -1.53125)        
    2483 => 207,          -- (100110.110011 | -25.203125)   => (110.01111 | -1.53125)        
    2484 => 207,          -- (100110.110100 | -25.1875)     => (110.01111 | -1.53125)        
    2485 => 207,          -- (100110.110101 | -25.171875)   => (110.01111 | -1.53125)        
    2486 => 207,          -- (100110.110110 | -25.15625)    => (110.01111 | -1.53125)        
    2487 => 207,          -- (100110.110111 | -25.140625)   => (110.01111 | -1.53125)        
    2488 => 207,          -- (100110.111000 | -25.125)      => (110.01111 | -1.53125)        
    2489 => 207,          -- (100110.111001 | -25.109375)   => (110.01111 | -1.53125)        
    2490 => 207,          -- (100110.111010 | -25.09375)    => (110.01111 | -1.53125)        
    2491 => 207,          -- (100110.111011 | -25.078125)   => (110.01111 | -1.53125)        
    2492 => 207,          -- (100110.111100 | -25.0625)     => (110.01111 | -1.53125)        
    2493 => 207,          -- (100110.111101 | -25.046875)   => (110.01111 | -1.53125)        
    2494 => 207,          -- (100110.111110 | -25.03125)    => (110.01111 | -1.53125)        
    2495 => 207,          -- (100110.111111 | -25.015625)   => (110.01111 | -1.53125)        
    2496 => 207,          -- (100111.000000 | -25.0)        => (110.01111 | -1.53125)        
    2497 => 207,          -- (100111.000001 | -24.984375)   => (110.01111 | -1.53125)        
    2498 => 207,          -- (100111.000010 | -24.96875)    => (110.01111 | -1.53125)        
    2499 => 207,          -- (100111.000011 | -24.953125)   => (110.01111 | -1.53125)        
    2500 => 207,          -- (100111.000100 | -24.9375)     => (110.01111 | -1.53125)        
    2501 => 207,          -- (100111.000101 | -24.921875)   => (110.01111 | -1.53125)        
    2502 => 207,          -- (100111.000110 | -24.90625)    => (110.01111 | -1.53125)        
    2503 => 207,          -- (100111.000111 | -24.890625)   => (110.01111 | -1.53125)        
    2504 => 207,          -- (100111.001000 | -24.875)      => (110.01111 | -1.53125)        
    2505 => 207,          -- (100111.001001 | -24.859375)   => (110.01111 | -1.53125)        
    2506 => 207,          -- (100111.001010 | -24.84375)    => (110.01111 | -1.53125)        
    2507 => 207,          -- (100111.001011 | -24.828125)   => (110.01111 | -1.53125)        
    2508 => 207,          -- (100111.001100 | -24.8125)     => (110.01111 | -1.53125)        
    2509 => 207,          -- (100111.001101 | -24.796875)   => (110.01111 | -1.53125)        
    2510 => 207,          -- (100111.001110 | -24.78125)    => (110.01111 | -1.53125)        
    2511 => 207,          -- (100111.001111 | -24.765625)   => (110.01111 | -1.53125)        
    2512 => 207,          -- (100111.010000 | -24.75)       => (110.01111 | -1.53125)        
    2513 => 207,          -- (100111.010001 | -24.734375)   => (110.01111 | -1.53125)        
    2514 => 207,          -- (100111.010010 | -24.71875)    => (110.01111 | -1.53125)        
    2515 => 207,          -- (100111.010011 | -24.703125)   => (110.01111 | -1.53125)        
    2516 => 207,          -- (100111.010100 | -24.6875)     => (110.01111 | -1.53125)        
    2517 => 207,          -- (100111.010101 | -24.671875)   => (110.01111 | -1.53125)        
    2518 => 207,          -- (100111.010110 | -24.65625)    => (110.01111 | -1.53125)        
    2519 => 207,          -- (100111.010111 | -24.640625)   => (110.01111 | -1.53125)        
    2520 => 207,          -- (100111.011000 | -24.625)      => (110.01111 | -1.53125)        
    2521 => 207,          -- (100111.011001 | -24.609375)   => (110.01111 | -1.53125)        
    2522 => 207,          -- (100111.011010 | -24.59375)    => (110.01111 | -1.53125)        
    2523 => 207,          -- (100111.011011 | -24.578125)   => (110.01111 | -1.53125)        
    2524 => 207,          -- (100111.011100 | -24.5625)     => (110.01111 | -1.53125)        
    2525 => 207,          -- (100111.011101 | -24.546875)   => (110.01111 | -1.53125)        
    2526 => 207,          -- (100111.011110 | -24.53125)    => (110.01111 | -1.53125)        
    2527 => 207,          -- (100111.011111 | -24.515625)   => (110.01111 | -1.53125)        
    2528 => 207,          -- (100111.100000 | -24.5)        => (110.01111 | -1.53125)        
    2529 => 207,          -- (100111.100001 | -24.484375)   => (110.01111 | -1.53125)        
    2530 => 207,          -- (100111.100010 | -24.46875)    => (110.01111 | -1.53125)        
    2531 => 207,          -- (100111.100011 | -24.453125)   => (110.01111 | -1.53125)        
    2532 => 207,          -- (100111.100100 | -24.4375)     => (110.01111 | -1.53125)        
    2533 => 207,          -- (100111.100101 | -24.421875)   => (110.01111 | -1.53125)        
    2534 => 207,          -- (100111.100110 | -24.40625)    => (110.01111 | -1.53125)        
    2535 => 207,          -- (100111.100111 | -24.390625)   => (110.01111 | -1.53125)        
    2536 => 207,          -- (100111.101000 | -24.375)      => (110.01111 | -1.53125)        
    2537 => 207,          -- (100111.101001 | -24.359375)   => (110.01111 | -1.53125)        
    2538 => 207,          -- (100111.101010 | -24.34375)    => (110.01111 | -1.53125)        
    2539 => 207,          -- (100111.101011 | -24.328125)   => (110.01111 | -1.53125)        
    2540 => 207,          -- (100111.101100 | -24.3125)     => (110.01111 | -1.53125)        
    2541 => 207,          -- (100111.101101 | -24.296875)   => (110.01111 | -1.53125)        
    2542 => 207,          -- (100111.101110 | -24.28125)    => (110.01111 | -1.53125)        
    2543 => 207,          -- (100111.101111 | -24.265625)   => (110.01111 | -1.53125)        
    2544 => 207,          -- (100111.110000 | -24.25)       => (110.01111 | -1.53125)        
    2545 => 207,          -- (100111.110001 | -24.234375)   => (110.01111 | -1.53125)        
    2546 => 207,          -- (100111.110010 | -24.21875)    => (110.01111 | -1.53125)        
    2547 => 207,          -- (100111.110011 | -24.203125)   => (110.01111 | -1.53125)        
    2548 => 207,          -- (100111.110100 | -24.1875)     => (110.01111 | -1.53125)        
    2549 => 207,          -- (100111.110101 | -24.171875)   => (110.01111 | -1.53125)        
    2550 => 207,          -- (100111.110110 | -24.15625)    => (110.01111 | -1.53125)        
    2551 => 207,          -- (100111.110111 | -24.140625)   => (110.01111 | -1.53125)        
    2552 => 207,          -- (100111.111000 | -24.125)      => (110.01111 | -1.53125)        
    2553 => 207,          -- (100111.111001 | -24.109375)   => (110.01111 | -1.53125)        
    2554 => 207,          -- (100111.111010 | -24.09375)    => (110.01111 | -1.53125)        
    2555 => 207,          -- (100111.111011 | -24.078125)   => (110.01111 | -1.53125)        
    2556 => 207,          -- (100111.111100 | -24.0625)     => (110.01111 | -1.53125)        
    2557 => 207,          -- (100111.111101 | -24.046875)   => (110.01111 | -1.53125)        
    2558 => 207,          -- (100111.111110 | -24.03125)    => (110.01111 | -1.53125)        
    2559 => 207,          -- (100111.111111 | -24.015625)   => (110.01111 | -1.53125)        
    2560 => 207,          -- (101000.000000 | -24.0)        => (110.01111 | -1.53125)        
    2561 => 207,          -- (101000.000001 | -23.984375)   => (110.01111 | -1.53125)        
    2562 => 207,          -- (101000.000010 | -23.96875)    => (110.01111 | -1.53125)        
    2563 => 207,          -- (101000.000011 | -23.953125)   => (110.01111 | -1.53125)        
    2564 => 207,          -- (101000.000100 | -23.9375)     => (110.01111 | -1.53125)        
    2565 => 207,          -- (101000.000101 | -23.921875)   => (110.01111 | -1.53125)        
    2566 => 207,          -- (101000.000110 | -23.90625)    => (110.01111 | -1.53125)        
    2567 => 207,          -- (101000.000111 | -23.890625)   => (110.01111 | -1.53125)        
    2568 => 207,          -- (101000.001000 | -23.875)      => (110.01111 | -1.53125)        
    2569 => 207,          -- (101000.001001 | -23.859375)   => (110.01111 | -1.53125)        
    2570 => 207,          -- (101000.001010 | -23.84375)    => (110.01111 | -1.53125)        
    2571 => 207,          -- (101000.001011 | -23.828125)   => (110.01111 | -1.53125)        
    2572 => 207,          -- (101000.001100 | -23.8125)     => (110.01111 | -1.53125)        
    2573 => 207,          -- (101000.001101 | -23.796875)   => (110.01111 | -1.53125)        
    2574 => 207,          -- (101000.001110 | -23.78125)    => (110.01111 | -1.53125)        
    2575 => 207,          -- (101000.001111 | -23.765625)   => (110.01111 | -1.53125)        
    2576 => 207,          -- (101000.010000 | -23.75)       => (110.01111 | -1.53125)        
    2577 => 207,          -- (101000.010001 | -23.734375)   => (110.01111 | -1.53125)        
    2578 => 207,          -- (101000.010010 | -23.71875)    => (110.01111 | -1.53125)        
    2579 => 207,          -- (101000.010011 | -23.703125)   => (110.01111 | -1.53125)        
    2580 => 207,          -- (101000.010100 | -23.6875)     => (110.01111 | -1.53125)        
    2581 => 207,          -- (101000.010101 | -23.671875)   => (110.01111 | -1.53125)        
    2582 => 207,          -- (101000.010110 | -23.65625)    => (110.01111 | -1.53125)        
    2583 => 207,          -- (101000.010111 | -23.640625)   => (110.01111 | -1.53125)        
    2584 => 207,          -- (101000.011000 | -23.625)      => (110.01111 | -1.53125)        
    2585 => 207,          -- (101000.011001 | -23.609375)   => (110.01111 | -1.53125)        
    2586 => 207,          -- (101000.011010 | -23.59375)    => (110.01111 | -1.53125)        
    2587 => 207,          -- (101000.011011 | -23.578125)   => (110.01111 | -1.53125)        
    2588 => 207,          -- (101000.011100 | -23.5625)     => (110.01111 | -1.53125)        
    2589 => 207,          -- (101000.011101 | -23.546875)   => (110.01111 | -1.53125)        
    2590 => 207,          -- (101000.011110 | -23.53125)    => (110.01111 | -1.53125)        
    2591 => 207,          -- (101000.011111 | -23.515625)   => (110.01111 | -1.53125)        
    2592 => 207,          -- (101000.100000 | -23.5)        => (110.01111 | -1.53125)        
    2593 => 207,          -- (101000.100001 | -23.484375)   => (110.01111 | -1.53125)        
    2594 => 207,          -- (101000.100010 | -23.46875)    => (110.01111 | -1.53125)        
    2595 => 207,          -- (101000.100011 | -23.453125)   => (110.01111 | -1.53125)        
    2596 => 207,          -- (101000.100100 | -23.4375)     => (110.01111 | -1.53125)        
    2597 => 207,          -- (101000.100101 | -23.421875)   => (110.01111 | -1.53125)        
    2598 => 207,          -- (101000.100110 | -23.40625)    => (110.01111 | -1.53125)        
    2599 => 207,          -- (101000.100111 | -23.390625)   => (110.01111 | -1.53125)        
    2600 => 207,          -- (101000.101000 | -23.375)      => (110.01111 | -1.53125)        
    2601 => 207,          -- (101000.101001 | -23.359375)   => (110.01111 | -1.53125)        
    2602 => 207,          -- (101000.101010 | -23.34375)    => (110.01111 | -1.53125)        
    2603 => 207,          -- (101000.101011 | -23.328125)   => (110.01111 | -1.53125)        
    2604 => 207,          -- (101000.101100 | -23.3125)     => (110.01111 | -1.53125)        
    2605 => 207,          -- (101000.101101 | -23.296875)   => (110.01111 | -1.53125)        
    2606 => 207,          -- (101000.101110 | -23.28125)    => (110.01111 | -1.53125)        
    2607 => 207,          -- (101000.101111 | -23.265625)   => (110.01111 | -1.53125)        
    2608 => 207,          -- (101000.110000 | -23.25)       => (110.01111 | -1.53125)        
    2609 => 207,          -- (101000.110001 | -23.234375)   => (110.01111 | -1.53125)        
    2610 => 207,          -- (101000.110010 | -23.21875)    => (110.01111 | -1.53125)        
    2611 => 207,          -- (101000.110011 | -23.203125)   => (110.01111 | -1.53125)        
    2612 => 207,          -- (101000.110100 | -23.1875)     => (110.01111 | -1.53125)        
    2613 => 207,          -- (101000.110101 | -23.171875)   => (110.01111 | -1.53125)        
    2614 => 207,          -- (101000.110110 | -23.15625)    => (110.01111 | -1.53125)        
    2615 => 207,          -- (101000.110111 | -23.140625)   => (110.01111 | -1.53125)        
    2616 => 207,          -- (101000.111000 | -23.125)      => (110.01111 | -1.53125)        
    2617 => 207,          -- (101000.111001 | -23.109375)   => (110.01111 | -1.53125)        
    2618 => 207,          -- (101000.111010 | -23.09375)    => (110.01111 | -1.53125)        
    2619 => 207,          -- (101000.111011 | -23.078125)   => (110.01111 | -1.53125)        
    2620 => 207,          -- (101000.111100 | -23.0625)     => (110.01111 | -1.53125)        
    2621 => 207,          -- (101000.111101 | -23.046875)   => (110.01111 | -1.53125)        
    2622 => 207,          -- (101000.111110 | -23.03125)    => (110.01111 | -1.53125)        
    2623 => 207,          -- (101000.111111 | -23.015625)   => (110.01111 | -1.53125)        
    2624 => 207,          -- (101001.000000 | -23.0)        => (110.01111 | -1.53125)        
    2625 => 207,          -- (101001.000001 | -22.984375)   => (110.01111 | -1.53125)        
    2626 => 207,          -- (101001.000010 | -22.96875)    => (110.01111 | -1.53125)        
    2627 => 207,          -- (101001.000011 | -22.953125)   => (110.01111 | -1.53125)        
    2628 => 207,          -- (101001.000100 | -22.9375)     => (110.01111 | -1.53125)        
    2629 => 207,          -- (101001.000101 | -22.921875)   => (110.01111 | -1.53125)        
    2630 => 207,          -- (101001.000110 | -22.90625)    => (110.01111 | -1.53125)        
    2631 => 207,          -- (101001.000111 | -22.890625)   => (110.01111 | -1.53125)        
    2632 => 207,          -- (101001.001000 | -22.875)      => (110.01111 | -1.53125)        
    2633 => 207,          -- (101001.001001 | -22.859375)   => (110.01111 | -1.53125)        
    2634 => 207,          -- (101001.001010 | -22.84375)    => (110.01111 | -1.53125)        
    2635 => 207,          -- (101001.001011 | -22.828125)   => (110.01111 | -1.53125)        
    2636 => 207,          -- (101001.001100 | -22.8125)     => (110.01111 | -1.53125)        
    2637 => 207,          -- (101001.001101 | -22.796875)   => (110.01111 | -1.53125)        
    2638 => 207,          -- (101001.001110 | -22.78125)    => (110.01111 | -1.53125)        
    2639 => 207,          -- (101001.001111 | -22.765625)   => (110.01111 | -1.53125)        
    2640 => 207,          -- (101001.010000 | -22.75)       => (110.01111 | -1.53125)        
    2641 => 207,          -- (101001.010001 | -22.734375)   => (110.01111 | -1.53125)        
    2642 => 207,          -- (101001.010010 | -22.71875)    => (110.01111 | -1.53125)        
    2643 => 207,          -- (101001.010011 | -22.703125)   => (110.01111 | -1.53125)        
    2644 => 207,          -- (101001.010100 | -22.6875)     => (110.01111 | -1.53125)        
    2645 => 207,          -- (101001.010101 | -22.671875)   => (110.01111 | -1.53125)        
    2646 => 207,          -- (101001.010110 | -22.65625)    => (110.01111 | -1.53125)        
    2647 => 207,          -- (101001.010111 | -22.640625)   => (110.01111 | -1.53125)        
    2648 => 207,          -- (101001.011000 | -22.625)      => (110.01111 | -1.53125)        
    2649 => 207,          -- (101001.011001 | -22.609375)   => (110.01111 | -1.53125)        
    2650 => 207,          -- (101001.011010 | -22.59375)    => (110.01111 | -1.53125)        
    2651 => 207,          -- (101001.011011 | -22.578125)   => (110.01111 | -1.53125)        
    2652 => 207,          -- (101001.011100 | -22.5625)     => (110.01111 | -1.53125)        
    2653 => 207,          -- (101001.011101 | -22.546875)   => (110.01111 | -1.53125)        
    2654 => 207,          -- (101001.011110 | -22.53125)    => (110.01111 | -1.53125)        
    2655 => 207,          -- (101001.011111 | -22.515625)   => (110.01111 | -1.53125)        
    2656 => 207,          -- (101001.100000 | -22.5)        => (110.01111 | -1.53125)        
    2657 => 207,          -- (101001.100001 | -22.484375)   => (110.01111 | -1.53125)        
    2658 => 207,          -- (101001.100010 | -22.46875)    => (110.01111 | -1.53125)        
    2659 => 207,          -- (101001.100011 | -22.453125)   => (110.01111 | -1.53125)        
    2660 => 207,          -- (101001.100100 | -22.4375)     => (110.01111 | -1.53125)        
    2661 => 207,          -- (101001.100101 | -22.421875)   => (110.01111 | -1.53125)        
    2662 => 207,          -- (101001.100110 | -22.40625)    => (110.01111 | -1.53125)        
    2663 => 207,          -- (101001.100111 | -22.390625)   => (110.01111 | -1.53125)        
    2664 => 207,          -- (101001.101000 | -22.375)      => (110.01111 | -1.53125)        
    2665 => 207,          -- (101001.101001 | -22.359375)   => (110.01111 | -1.53125)        
    2666 => 207,          -- (101001.101010 | -22.34375)    => (110.01111 | -1.53125)        
    2667 => 207,          -- (101001.101011 | -22.328125)   => (110.01111 | -1.53125)        
    2668 => 207,          -- (101001.101100 | -22.3125)     => (110.01111 | -1.53125)        
    2669 => 207,          -- (101001.101101 | -22.296875)   => (110.01111 | -1.53125)        
    2670 => 207,          -- (101001.101110 | -22.28125)    => (110.01111 | -1.53125)        
    2671 => 207,          -- (101001.101111 | -22.265625)   => (110.01111 | -1.53125)        
    2672 => 207,          -- (101001.110000 | -22.25)       => (110.01111 | -1.53125)        
    2673 => 207,          -- (101001.110001 | -22.234375)   => (110.01111 | -1.53125)        
    2674 => 207,          -- (101001.110010 | -22.21875)    => (110.01111 | -1.53125)        
    2675 => 207,          -- (101001.110011 | -22.203125)   => (110.01111 | -1.53125)        
    2676 => 207,          -- (101001.110100 | -22.1875)     => (110.01111 | -1.53125)        
    2677 => 207,          -- (101001.110101 | -22.171875)   => (110.01111 | -1.53125)        
    2678 => 207,          -- (101001.110110 | -22.15625)    => (110.01111 | -1.53125)        
    2679 => 207,          -- (101001.110111 | -22.140625)   => (110.01111 | -1.53125)        
    2680 => 207,          -- (101001.111000 | -22.125)      => (110.01111 | -1.53125)        
    2681 => 207,          -- (101001.111001 | -22.109375)   => (110.01111 | -1.53125)        
    2682 => 207,          -- (101001.111010 | -22.09375)    => (110.01111 | -1.53125)        
    2683 => 207,          -- (101001.111011 | -22.078125)   => (110.01111 | -1.53125)        
    2684 => 207,          -- (101001.111100 | -22.0625)     => (110.01111 | -1.53125)        
    2685 => 207,          -- (101001.111101 | -22.046875)   => (110.01111 | -1.53125)        
    2686 => 207,          -- (101001.111110 | -22.03125)    => (110.01111 | -1.53125)        
    2687 => 207,          -- (101001.111111 | -22.015625)   => (110.01111 | -1.53125)        
    2688 => 207,          -- (101010.000000 | -22.0)        => (110.01111 | -1.53125)        
    2689 => 207,          -- (101010.000001 | -21.984375)   => (110.01111 | -1.53125)        
    2690 => 207,          -- (101010.000010 | -21.96875)    => (110.01111 | -1.53125)        
    2691 => 207,          -- (101010.000011 | -21.953125)   => (110.01111 | -1.53125)        
    2692 => 207,          -- (101010.000100 | -21.9375)     => (110.01111 | -1.53125)        
    2693 => 207,          -- (101010.000101 | -21.921875)   => (110.01111 | -1.53125)        
    2694 => 207,          -- (101010.000110 | -21.90625)    => (110.01111 | -1.53125)        
    2695 => 207,          -- (101010.000111 | -21.890625)   => (110.01111 | -1.53125)        
    2696 => 207,          -- (101010.001000 | -21.875)      => (110.01111 | -1.53125)        
    2697 => 207,          -- (101010.001001 | -21.859375)   => (110.01111 | -1.53125)        
    2698 => 207,          -- (101010.001010 | -21.84375)    => (110.01111 | -1.53125)        
    2699 => 207,          -- (101010.001011 | -21.828125)   => (110.01111 | -1.53125)        
    2700 => 207,          -- (101010.001100 | -21.8125)     => (110.01111 | -1.53125)        
    2701 => 207,          -- (101010.001101 | -21.796875)   => (110.01111 | -1.53125)        
    2702 => 207,          -- (101010.001110 | -21.78125)    => (110.01111 | -1.53125)        
    2703 => 207,          -- (101010.001111 | -21.765625)   => (110.01111 | -1.53125)        
    2704 => 207,          -- (101010.010000 | -21.75)       => (110.01111 | -1.53125)        
    2705 => 207,          -- (101010.010001 | -21.734375)   => (110.01111 | -1.53125)        
    2706 => 207,          -- (101010.010010 | -21.71875)    => (110.01111 | -1.53125)        
    2707 => 207,          -- (101010.010011 | -21.703125)   => (110.01111 | -1.53125)        
    2708 => 207,          -- (101010.010100 | -21.6875)     => (110.01111 | -1.53125)        
    2709 => 207,          -- (101010.010101 | -21.671875)   => (110.01111 | -1.53125)        
    2710 => 207,          -- (101010.010110 | -21.65625)    => (110.01111 | -1.53125)        
    2711 => 207,          -- (101010.010111 | -21.640625)   => (110.01111 | -1.53125)        
    2712 => 207,          -- (101010.011000 | -21.625)      => (110.01111 | -1.53125)        
    2713 => 207,          -- (101010.011001 | -21.609375)   => (110.01111 | -1.53125)        
    2714 => 207,          -- (101010.011010 | -21.59375)    => (110.01111 | -1.53125)        
    2715 => 207,          -- (101010.011011 | -21.578125)   => (110.01111 | -1.53125)        
    2716 => 207,          -- (101010.011100 | -21.5625)     => (110.01111 | -1.53125)        
    2717 => 207,          -- (101010.011101 | -21.546875)   => (110.01111 | -1.53125)        
    2718 => 207,          -- (101010.011110 | -21.53125)    => (110.01111 | -1.53125)        
    2719 => 207,          -- (101010.011111 | -21.515625)   => (110.01111 | -1.53125)        
    2720 => 207,          -- (101010.100000 | -21.5)        => (110.01111 | -1.53125)        
    2721 => 207,          -- (101010.100001 | -21.484375)   => (110.01111 | -1.53125)        
    2722 => 207,          -- (101010.100010 | -21.46875)    => (110.01111 | -1.53125)        
    2723 => 207,          -- (101010.100011 | -21.453125)   => (110.01111 | -1.53125)        
    2724 => 207,          -- (101010.100100 | -21.4375)     => (110.01111 | -1.53125)        
    2725 => 207,          -- (101010.100101 | -21.421875)   => (110.01111 | -1.53125)        
    2726 => 207,          -- (101010.100110 | -21.40625)    => (110.01111 | -1.53125)        
    2727 => 207,          -- (101010.100111 | -21.390625)   => (110.01111 | -1.53125)        
    2728 => 207,          -- (101010.101000 | -21.375)      => (110.01111 | -1.53125)        
    2729 => 207,          -- (101010.101001 | -21.359375)   => (110.01111 | -1.53125)        
    2730 => 207,          -- (101010.101010 | -21.34375)    => (110.01111 | -1.53125)        
    2731 => 207,          -- (101010.101011 | -21.328125)   => (110.01111 | -1.53125)        
    2732 => 207,          -- (101010.101100 | -21.3125)     => (110.01111 | -1.53125)        
    2733 => 207,          -- (101010.101101 | -21.296875)   => (110.01111 | -1.53125)        
    2734 => 207,          -- (101010.101110 | -21.28125)    => (110.01111 | -1.53125)        
    2735 => 207,          -- (101010.101111 | -21.265625)   => (110.01111 | -1.53125)        
    2736 => 207,          -- (101010.110000 | -21.25)       => (110.01111 | -1.53125)        
    2737 => 207,          -- (101010.110001 | -21.234375)   => (110.01111 | -1.53125)        
    2738 => 207,          -- (101010.110010 | -21.21875)    => (110.01111 | -1.53125)        
    2739 => 207,          -- (101010.110011 | -21.203125)   => (110.01111 | -1.53125)        
    2740 => 207,          -- (101010.110100 | -21.1875)     => (110.01111 | -1.53125)        
    2741 => 207,          -- (101010.110101 | -21.171875)   => (110.01111 | -1.53125)        
    2742 => 207,          -- (101010.110110 | -21.15625)    => (110.01111 | -1.53125)        
    2743 => 207,          -- (101010.110111 | -21.140625)   => (110.01111 | -1.53125)        
    2744 => 207,          -- (101010.111000 | -21.125)      => (110.01111 | -1.53125)        
    2745 => 207,          -- (101010.111001 | -21.109375)   => (110.01111 | -1.53125)        
    2746 => 207,          -- (101010.111010 | -21.09375)    => (110.01111 | -1.53125)        
    2747 => 207,          -- (101010.111011 | -21.078125)   => (110.01111 | -1.53125)        
    2748 => 207,          -- (101010.111100 | -21.0625)     => (110.01111 | -1.53125)        
    2749 => 207,          -- (101010.111101 | -21.046875)   => (110.01111 | -1.53125)        
    2750 => 207,          -- (101010.111110 | -21.03125)    => (110.01111 | -1.53125)        
    2751 => 207,          -- (101010.111111 | -21.015625)   => (110.01111 | -1.53125)        
    2752 => 207,          -- (101011.000000 | -21.0)        => (110.01111 | -1.53125)        
    2753 => 207,          -- (101011.000001 | -20.984375)   => (110.01111 | -1.53125)        
    2754 => 207,          -- (101011.000010 | -20.96875)    => (110.01111 | -1.53125)        
    2755 => 207,          -- (101011.000011 | -20.953125)   => (110.01111 | -1.53125)        
    2756 => 207,          -- (101011.000100 | -20.9375)     => (110.01111 | -1.53125)        
    2757 => 207,          -- (101011.000101 | -20.921875)   => (110.01111 | -1.53125)        
    2758 => 207,          -- (101011.000110 | -20.90625)    => (110.01111 | -1.53125)        
    2759 => 207,          -- (101011.000111 | -20.890625)   => (110.01111 | -1.53125)        
    2760 => 207,          -- (101011.001000 | -20.875)      => (110.01111 | -1.53125)        
    2761 => 207,          -- (101011.001001 | -20.859375)   => (110.01111 | -1.53125)        
    2762 => 207,          -- (101011.001010 | -20.84375)    => (110.01111 | -1.53125)        
    2763 => 207,          -- (101011.001011 | -20.828125)   => (110.01111 | -1.53125)        
    2764 => 207,          -- (101011.001100 | -20.8125)     => (110.01111 | -1.53125)        
    2765 => 207,          -- (101011.001101 | -20.796875)   => (110.01111 | -1.53125)        
    2766 => 207,          -- (101011.001110 | -20.78125)    => (110.01111 | -1.53125)        
    2767 => 207,          -- (101011.001111 | -20.765625)   => (110.01111 | -1.53125)        
    2768 => 207,          -- (101011.010000 | -20.75)       => (110.01111 | -1.53125)        
    2769 => 207,          -- (101011.010001 | -20.734375)   => (110.01111 | -1.53125)        
    2770 => 207,          -- (101011.010010 | -20.71875)    => (110.01111 | -1.53125)        
    2771 => 207,          -- (101011.010011 | -20.703125)   => (110.01111 | -1.53125)        
    2772 => 207,          -- (101011.010100 | -20.6875)     => (110.01111 | -1.53125)        
    2773 => 207,          -- (101011.010101 | -20.671875)   => (110.01111 | -1.53125)        
    2774 => 207,          -- (101011.010110 | -20.65625)    => (110.01111 | -1.53125)        
    2775 => 207,          -- (101011.010111 | -20.640625)   => (110.01111 | -1.53125)        
    2776 => 207,          -- (101011.011000 | -20.625)      => (110.01111 | -1.53125)        
    2777 => 207,          -- (101011.011001 | -20.609375)   => (110.01111 | -1.53125)        
    2778 => 207,          -- (101011.011010 | -20.59375)    => (110.01111 | -1.53125)        
    2779 => 207,          -- (101011.011011 | -20.578125)   => (110.01111 | -1.53125)        
    2780 => 207,          -- (101011.011100 | -20.5625)     => (110.01111 | -1.53125)        
    2781 => 207,          -- (101011.011101 | -20.546875)   => (110.01111 | -1.53125)        
    2782 => 207,          -- (101011.011110 | -20.53125)    => (110.01111 | -1.53125)        
    2783 => 207,          -- (101011.011111 | -20.515625)   => (110.01111 | -1.53125)        
    2784 => 207,          -- (101011.100000 | -20.5)        => (110.01111 | -1.53125)        
    2785 => 207,          -- (101011.100001 | -20.484375)   => (110.01111 | -1.53125)        
    2786 => 207,          -- (101011.100010 | -20.46875)    => (110.01111 | -1.53125)        
    2787 => 207,          -- (101011.100011 | -20.453125)   => (110.01111 | -1.53125)        
    2788 => 207,          -- (101011.100100 | -20.4375)     => (110.01111 | -1.53125)        
    2789 => 207,          -- (101011.100101 | -20.421875)   => (110.01111 | -1.53125)        
    2790 => 207,          -- (101011.100110 | -20.40625)    => (110.01111 | -1.53125)        
    2791 => 207,          -- (101011.100111 | -20.390625)   => (110.01111 | -1.53125)        
    2792 => 207,          -- (101011.101000 | -20.375)      => (110.01111 | -1.53125)        
    2793 => 207,          -- (101011.101001 | -20.359375)   => (110.01111 | -1.53125)        
    2794 => 207,          -- (101011.101010 | -20.34375)    => (110.01111 | -1.53125)        
    2795 => 207,          -- (101011.101011 | -20.328125)   => (110.01111 | -1.53125)        
    2796 => 207,          -- (101011.101100 | -20.3125)     => (110.01111 | -1.53125)        
    2797 => 207,          -- (101011.101101 | -20.296875)   => (110.01111 | -1.53125)        
    2798 => 207,          -- (101011.101110 | -20.28125)    => (110.01111 | -1.53125)        
    2799 => 207,          -- (101011.101111 | -20.265625)   => (110.01111 | -1.53125)        
    2800 => 207,          -- (101011.110000 | -20.25)       => (110.01111 | -1.53125)        
    2801 => 207,          -- (101011.110001 | -20.234375)   => (110.01111 | -1.53125)        
    2802 => 207,          -- (101011.110010 | -20.21875)    => (110.01111 | -1.53125)        
    2803 => 207,          -- (101011.110011 | -20.203125)   => (110.01111 | -1.53125)        
    2804 => 207,          -- (101011.110100 | -20.1875)     => (110.01111 | -1.53125)        
    2805 => 207,          -- (101011.110101 | -20.171875)   => (110.01111 | -1.53125)        
    2806 => 207,          -- (101011.110110 | -20.15625)    => (110.01111 | -1.53125)        
    2807 => 207,          -- (101011.110111 | -20.140625)   => (110.01111 | -1.53125)        
    2808 => 207,          -- (101011.111000 | -20.125)      => (110.01111 | -1.53125)        
    2809 => 207,          -- (101011.111001 | -20.109375)   => (110.01111 | -1.53125)        
    2810 => 207,          -- (101011.111010 | -20.09375)    => (110.01111 | -1.53125)        
    2811 => 207,          -- (101011.111011 | -20.078125)   => (110.01111 | -1.53125)        
    2812 => 207,          -- (101011.111100 | -20.0625)     => (110.01111 | -1.53125)        
    2813 => 207,          -- (101011.111101 | -20.046875)   => (110.01111 | -1.53125)        
    2814 => 207,          -- (101011.111110 | -20.03125)    => (110.01111 | -1.53125)        
    2815 => 207,          -- (101011.111111 | -20.015625)   => (110.01111 | -1.53125)        
    2816 => 207,          -- (101100.000000 | -20.0)        => (110.01111 | -1.53125)        
    2817 => 207,          -- (101100.000001 | -19.984375)   => (110.01111 | -1.53125)        
    2818 => 207,          -- (101100.000010 | -19.96875)    => (110.01111 | -1.53125)        
    2819 => 207,          -- (101100.000011 | -19.953125)   => (110.01111 | -1.53125)        
    2820 => 207,          -- (101100.000100 | -19.9375)     => (110.01111 | -1.53125)        
    2821 => 207,          -- (101100.000101 | -19.921875)   => (110.01111 | -1.53125)        
    2822 => 207,          -- (101100.000110 | -19.90625)    => (110.01111 | -1.53125)        
    2823 => 207,          -- (101100.000111 | -19.890625)   => (110.01111 | -1.53125)        
    2824 => 207,          -- (101100.001000 | -19.875)      => (110.01111 | -1.53125)        
    2825 => 207,          -- (101100.001001 | -19.859375)   => (110.01111 | -1.53125)        
    2826 => 207,          -- (101100.001010 | -19.84375)    => (110.01111 | -1.53125)        
    2827 => 207,          -- (101100.001011 | -19.828125)   => (110.01111 | -1.53125)        
    2828 => 207,          -- (101100.001100 | -19.8125)     => (110.01111 | -1.53125)        
    2829 => 207,          -- (101100.001101 | -19.796875)   => (110.01111 | -1.53125)        
    2830 => 207,          -- (101100.001110 | -19.78125)    => (110.01111 | -1.53125)        
    2831 => 207,          -- (101100.001111 | -19.765625)   => (110.01111 | -1.53125)        
    2832 => 207,          -- (101100.010000 | -19.75)       => (110.01111 | -1.53125)        
    2833 => 207,          -- (101100.010001 | -19.734375)   => (110.01111 | -1.53125)        
    2834 => 207,          -- (101100.010010 | -19.71875)    => (110.01111 | -1.53125)        
    2835 => 207,          -- (101100.010011 | -19.703125)   => (110.01111 | -1.53125)        
    2836 => 207,          -- (101100.010100 | -19.6875)     => (110.01111 | -1.53125)        
    2837 => 207,          -- (101100.010101 | -19.671875)   => (110.01111 | -1.53125)        
    2838 => 207,          -- (101100.010110 | -19.65625)    => (110.01111 | -1.53125)        
    2839 => 207,          -- (101100.010111 | -19.640625)   => (110.01111 | -1.53125)        
    2840 => 207,          -- (101100.011000 | -19.625)      => (110.01111 | -1.53125)        
    2841 => 207,          -- (101100.011001 | -19.609375)   => (110.01111 | -1.53125)        
    2842 => 207,          -- (101100.011010 | -19.59375)    => (110.01111 | -1.53125)        
    2843 => 207,          -- (101100.011011 | -19.578125)   => (110.01111 | -1.53125)        
    2844 => 207,          -- (101100.011100 | -19.5625)     => (110.01111 | -1.53125)        
    2845 => 207,          -- (101100.011101 | -19.546875)   => (110.01111 | -1.53125)        
    2846 => 207,          -- (101100.011110 | -19.53125)    => (110.01111 | -1.53125)        
    2847 => 207,          -- (101100.011111 | -19.515625)   => (110.01111 | -1.53125)        
    2848 => 207,          -- (101100.100000 | -19.5)        => (110.01111 | -1.53125)        
    2849 => 207,          -- (101100.100001 | -19.484375)   => (110.01111 | -1.53125)        
    2850 => 207,          -- (101100.100010 | -19.46875)    => (110.01111 | -1.53125)        
    2851 => 207,          -- (101100.100011 | -19.453125)   => (110.01111 | -1.53125)        
    2852 => 207,          -- (101100.100100 | -19.4375)     => (110.01111 | -1.53125)        
    2853 => 207,          -- (101100.100101 | -19.421875)   => (110.01111 | -1.53125)        
    2854 => 207,          -- (101100.100110 | -19.40625)    => (110.01111 | -1.53125)        
    2855 => 207,          -- (101100.100111 | -19.390625)   => (110.01111 | -1.53125)        
    2856 => 207,          -- (101100.101000 | -19.375)      => (110.01111 | -1.53125)        
    2857 => 207,          -- (101100.101001 | -19.359375)   => (110.01111 | -1.53125)        
    2858 => 207,          -- (101100.101010 | -19.34375)    => (110.01111 | -1.53125)        
    2859 => 207,          -- (101100.101011 | -19.328125)   => (110.01111 | -1.53125)        
    2860 => 207,          -- (101100.101100 | -19.3125)     => (110.01111 | -1.53125)        
    2861 => 207,          -- (101100.101101 | -19.296875)   => (110.01111 | -1.53125)        
    2862 => 207,          -- (101100.101110 | -19.28125)    => (110.01111 | -1.53125)        
    2863 => 207,          -- (101100.101111 | -19.265625)   => (110.01111 | -1.53125)        
    2864 => 207,          -- (101100.110000 | -19.25)       => (110.01111 | -1.53125)        
    2865 => 207,          -- (101100.110001 | -19.234375)   => (110.01111 | -1.53125)        
    2866 => 207,          -- (101100.110010 | -19.21875)    => (110.01111 | -1.53125)        
    2867 => 207,          -- (101100.110011 | -19.203125)   => (110.01111 | -1.53125)        
    2868 => 207,          -- (101100.110100 | -19.1875)     => (110.01111 | -1.53125)        
    2869 => 207,          -- (101100.110101 | -19.171875)   => (110.01111 | -1.53125)        
    2870 => 207,          -- (101100.110110 | -19.15625)    => (110.01111 | -1.53125)        
    2871 => 207,          -- (101100.110111 | -19.140625)   => (110.01111 | -1.53125)        
    2872 => 207,          -- (101100.111000 | -19.125)      => (110.01111 | -1.53125)        
    2873 => 207,          -- (101100.111001 | -19.109375)   => (110.01111 | -1.53125)        
    2874 => 207,          -- (101100.111010 | -19.09375)    => (110.01111 | -1.53125)        
    2875 => 207,          -- (101100.111011 | -19.078125)   => (110.01111 | -1.53125)        
    2876 => 207,          -- (101100.111100 | -19.0625)     => (110.01111 | -1.53125)        
    2877 => 207,          -- (101100.111101 | -19.046875)   => (110.01111 | -1.53125)        
    2878 => 207,          -- (101100.111110 | -19.03125)    => (110.01111 | -1.53125)        
    2879 => 207,          -- (101100.111111 | -19.015625)   => (110.01111 | -1.53125)        
    2880 => 207,          -- (101101.000000 | -19.0)        => (110.01111 | -1.53125)        
    2881 => 207,          -- (101101.000001 | -18.984375)   => (110.01111 | -1.53125)        
    2882 => 207,          -- (101101.000010 | -18.96875)    => (110.01111 | -1.53125)        
    2883 => 207,          -- (101101.000011 | -18.953125)   => (110.01111 | -1.53125)        
    2884 => 207,          -- (101101.000100 | -18.9375)     => (110.01111 | -1.53125)        
    2885 => 207,          -- (101101.000101 | -18.921875)   => (110.01111 | -1.53125)        
    2886 => 207,          -- (101101.000110 | -18.90625)    => (110.01111 | -1.53125)        
    2887 => 207,          -- (101101.000111 | -18.890625)   => (110.01111 | -1.53125)        
    2888 => 207,          -- (101101.001000 | -18.875)      => (110.01111 | -1.53125)        
    2889 => 207,          -- (101101.001001 | -18.859375)   => (110.01111 | -1.53125)        
    2890 => 207,          -- (101101.001010 | -18.84375)    => (110.01111 | -1.53125)        
    2891 => 207,          -- (101101.001011 | -18.828125)   => (110.01111 | -1.53125)        
    2892 => 207,          -- (101101.001100 | -18.8125)     => (110.01111 | -1.53125)        
    2893 => 207,          -- (101101.001101 | -18.796875)   => (110.01111 | -1.53125)        
    2894 => 207,          -- (101101.001110 | -18.78125)    => (110.01111 | -1.53125)        
    2895 => 207,          -- (101101.001111 | -18.765625)   => (110.01111 | -1.53125)        
    2896 => 207,          -- (101101.010000 | -18.75)       => (110.01111 | -1.53125)        
    2897 => 207,          -- (101101.010001 | -18.734375)   => (110.01111 | -1.53125)        
    2898 => 207,          -- (101101.010010 | -18.71875)    => (110.01111 | -1.53125)        
    2899 => 207,          -- (101101.010011 | -18.703125)   => (110.01111 | -1.53125)        
    2900 => 207,          -- (101101.010100 | -18.6875)     => (110.01111 | -1.53125)        
    2901 => 207,          -- (101101.010101 | -18.671875)   => (110.01111 | -1.53125)        
    2902 => 207,          -- (101101.010110 | -18.65625)    => (110.01111 | -1.53125)        
    2903 => 207,          -- (101101.010111 | -18.640625)   => (110.01111 | -1.53125)        
    2904 => 207,          -- (101101.011000 | -18.625)      => (110.01111 | -1.53125)        
    2905 => 207,          -- (101101.011001 | -18.609375)   => (110.01111 | -1.53125)        
    2906 => 207,          -- (101101.011010 | -18.59375)    => (110.01111 | -1.53125)        
    2907 => 207,          -- (101101.011011 | -18.578125)   => (110.01111 | -1.53125)        
    2908 => 207,          -- (101101.011100 | -18.5625)     => (110.01111 | -1.53125)        
    2909 => 207,          -- (101101.011101 | -18.546875)   => (110.01111 | -1.53125)        
    2910 => 207,          -- (101101.011110 | -18.53125)    => (110.01111 | -1.53125)        
    2911 => 207,          -- (101101.011111 | -18.515625)   => (110.01111 | -1.53125)        
    2912 => 207,          -- (101101.100000 | -18.5)        => (110.01111 | -1.53125)        
    2913 => 207,          -- (101101.100001 | -18.484375)   => (110.01111 | -1.53125)        
    2914 => 207,          -- (101101.100010 | -18.46875)    => (110.01111 | -1.53125)        
    2915 => 207,          -- (101101.100011 | -18.453125)   => (110.01111 | -1.53125)        
    2916 => 207,          -- (101101.100100 | -18.4375)     => (110.01111 | -1.53125)        
    2917 => 207,          -- (101101.100101 | -18.421875)   => (110.01111 | -1.53125)        
    2918 => 207,          -- (101101.100110 | -18.40625)    => (110.01111 | -1.53125)        
    2919 => 207,          -- (101101.100111 | -18.390625)   => (110.01111 | -1.53125)        
    2920 => 207,          -- (101101.101000 | -18.375)      => (110.01111 | -1.53125)        
    2921 => 207,          -- (101101.101001 | -18.359375)   => (110.01111 | -1.53125)        
    2922 => 207,          -- (101101.101010 | -18.34375)    => (110.01111 | -1.53125)        
    2923 => 207,          -- (101101.101011 | -18.328125)   => (110.01111 | -1.53125)        
    2924 => 207,          -- (101101.101100 | -18.3125)     => (110.01111 | -1.53125)        
    2925 => 207,          -- (101101.101101 | -18.296875)   => (110.01111 | -1.53125)        
    2926 => 207,          -- (101101.101110 | -18.28125)    => (110.01111 | -1.53125)        
    2927 => 207,          -- (101101.101111 | -18.265625)   => (110.01111 | -1.53125)        
    2928 => 207,          -- (101101.110000 | -18.25)       => (110.01111 | -1.53125)        
    2929 => 207,          -- (101101.110001 | -18.234375)   => (110.01111 | -1.53125)        
    2930 => 207,          -- (101101.110010 | -18.21875)    => (110.01111 | -1.53125)        
    2931 => 207,          -- (101101.110011 | -18.203125)   => (110.01111 | -1.53125)        
    2932 => 207,          -- (101101.110100 | -18.1875)     => (110.01111 | -1.53125)        
    2933 => 207,          -- (101101.110101 | -18.171875)   => (110.01111 | -1.53125)        
    2934 => 207,          -- (101101.110110 | -18.15625)    => (110.01111 | -1.53125)        
    2935 => 207,          -- (101101.110111 | -18.140625)   => (110.01111 | -1.53125)        
    2936 => 207,          -- (101101.111000 | -18.125)      => (110.01111 | -1.53125)        
    2937 => 207,          -- (101101.111001 | -18.109375)   => (110.01111 | -1.53125)        
    2938 => 207,          -- (101101.111010 | -18.09375)    => (110.01111 | -1.53125)        
    2939 => 207,          -- (101101.111011 | -18.078125)   => (110.01111 | -1.53125)        
    2940 => 207,          -- (101101.111100 | -18.0625)     => (110.01111 | -1.53125)        
    2941 => 207,          -- (101101.111101 | -18.046875)   => (110.01111 | -1.53125)        
    2942 => 207,          -- (101101.111110 | -18.03125)    => (110.01111 | -1.53125)        
    2943 => 207,          -- (101101.111111 | -18.015625)   => (110.01111 | -1.53125)        
    2944 => 207,          -- (101110.000000 | -18.0)        => (110.01111 | -1.53125)        
    2945 => 207,          -- (101110.000001 | -17.984375)   => (110.01111 | -1.53125)        
    2946 => 207,          -- (101110.000010 | -17.96875)    => (110.01111 | -1.53125)        
    2947 => 207,          -- (101110.000011 | -17.953125)   => (110.01111 | -1.53125)        
    2948 => 207,          -- (101110.000100 | -17.9375)     => (110.01111 | -1.53125)        
    2949 => 207,          -- (101110.000101 | -17.921875)   => (110.01111 | -1.53125)        
    2950 => 207,          -- (101110.000110 | -17.90625)    => (110.01111 | -1.53125)        
    2951 => 207,          -- (101110.000111 | -17.890625)   => (110.01111 | -1.53125)        
    2952 => 207,          -- (101110.001000 | -17.875)      => (110.01111 | -1.53125)        
    2953 => 207,          -- (101110.001001 | -17.859375)   => (110.01111 | -1.53125)        
    2954 => 207,          -- (101110.001010 | -17.84375)    => (110.01111 | -1.53125)        
    2955 => 207,          -- (101110.001011 | -17.828125)   => (110.01111 | -1.53125)        
    2956 => 207,          -- (101110.001100 | -17.8125)     => (110.01111 | -1.53125)        
    2957 => 207,          -- (101110.001101 | -17.796875)   => (110.01111 | -1.53125)        
    2958 => 207,          -- (101110.001110 | -17.78125)    => (110.01111 | -1.53125)        
    2959 => 207,          -- (101110.001111 | -17.765625)   => (110.01111 | -1.53125)        
    2960 => 207,          -- (101110.010000 | -17.75)       => (110.01111 | -1.53125)        
    2961 => 207,          -- (101110.010001 | -17.734375)   => (110.01111 | -1.53125)        
    2962 => 207,          -- (101110.010010 | -17.71875)    => (110.01111 | -1.53125)        
    2963 => 207,          -- (101110.010011 | -17.703125)   => (110.01111 | -1.53125)        
    2964 => 207,          -- (101110.010100 | -17.6875)     => (110.01111 | -1.53125)        
    2965 => 207,          -- (101110.010101 | -17.671875)   => (110.01111 | -1.53125)        
    2966 => 207,          -- (101110.010110 | -17.65625)    => (110.01111 | -1.53125)        
    2967 => 207,          -- (101110.010111 | -17.640625)   => (110.01111 | -1.53125)        
    2968 => 207,          -- (101110.011000 | -17.625)      => (110.01111 | -1.53125)        
    2969 => 207,          -- (101110.011001 | -17.609375)   => (110.01111 | -1.53125)        
    2970 => 207,          -- (101110.011010 | -17.59375)    => (110.01111 | -1.53125)        
    2971 => 207,          -- (101110.011011 | -17.578125)   => (110.01111 | -1.53125)        
    2972 => 207,          -- (101110.011100 | -17.5625)     => (110.01111 | -1.53125)        
    2973 => 207,          -- (101110.011101 | -17.546875)   => (110.01111 | -1.53125)        
    2974 => 207,          -- (101110.011110 | -17.53125)    => (110.01111 | -1.53125)        
    2975 => 207,          -- (101110.011111 | -17.515625)   => (110.01111 | -1.53125)        
    2976 => 207,          -- (101110.100000 | -17.5)        => (110.01111 | -1.53125)        
    2977 => 207,          -- (101110.100001 | -17.484375)   => (110.01111 | -1.53125)        
    2978 => 207,          -- (101110.100010 | -17.46875)    => (110.01111 | -1.53125)        
    2979 => 207,          -- (101110.100011 | -17.453125)   => (110.01111 | -1.53125)        
    2980 => 207,          -- (101110.100100 | -17.4375)     => (110.01111 | -1.53125)        
    2981 => 207,          -- (101110.100101 | -17.421875)   => (110.01111 | -1.53125)        
    2982 => 207,          -- (101110.100110 | -17.40625)    => (110.01111 | -1.53125)        
    2983 => 207,          -- (101110.100111 | -17.390625)   => (110.01111 | -1.53125)        
    2984 => 207,          -- (101110.101000 | -17.375)      => (110.01111 | -1.53125)        
    2985 => 207,          -- (101110.101001 | -17.359375)   => (110.01111 | -1.53125)        
    2986 => 207,          -- (101110.101010 | -17.34375)    => (110.01111 | -1.53125)        
    2987 => 207,          -- (101110.101011 | -17.328125)   => (110.01111 | -1.53125)        
    2988 => 207,          -- (101110.101100 | -17.3125)     => (110.01111 | -1.53125)        
    2989 => 207,          -- (101110.101101 | -17.296875)   => (110.01111 | -1.53125)        
    2990 => 207,          -- (101110.101110 | -17.28125)    => (110.01111 | -1.53125)        
    2991 => 207,          -- (101110.101111 | -17.265625)   => (110.01111 | -1.53125)        
    2992 => 207,          -- (101110.110000 | -17.25)       => (110.01111 | -1.53125)        
    2993 => 207,          -- (101110.110001 | -17.234375)   => (110.01111 | -1.53125)        
    2994 => 207,          -- (101110.110010 | -17.21875)    => (110.01111 | -1.53125)        
    2995 => 207,          -- (101110.110011 | -17.203125)   => (110.01111 | -1.53125)        
    2996 => 207,          -- (101110.110100 | -17.1875)     => (110.01111 | -1.53125)        
    2997 => 207,          -- (101110.110101 | -17.171875)   => (110.01111 | -1.53125)        
    2998 => 207,          -- (101110.110110 | -17.15625)    => (110.01111 | -1.53125)        
    2999 => 207,          -- (101110.110111 | -17.140625)   => (110.01111 | -1.53125)        
    3000 => 207,          -- (101110.111000 | -17.125)      => (110.01111 | -1.53125)        
    3001 => 207,          -- (101110.111001 | -17.109375)   => (110.01111 | -1.53125)        
    3002 => 207,          -- (101110.111010 | -17.09375)    => (110.01111 | -1.53125)        
    3003 => 207,          -- (101110.111011 | -17.078125)   => (110.01111 | -1.53125)        
    3004 => 207,          -- (101110.111100 | -17.0625)     => (110.01111 | -1.53125)        
    3005 => 207,          -- (101110.111101 | -17.046875)   => (110.01111 | -1.53125)        
    3006 => 207,          -- (101110.111110 | -17.03125)    => (110.01111 | -1.53125)        
    3007 => 207,          -- (101110.111111 | -17.015625)   => (110.01111 | -1.53125)        
    3008 => 207,          -- (101111.000000 | -17.0)        => (110.01111 | -1.53125)        
    3009 => 207,          -- (101111.000001 | -16.984375)   => (110.01111 | -1.53125)        
    3010 => 207,          -- (101111.000010 | -16.96875)    => (110.01111 | -1.53125)        
    3011 => 207,          -- (101111.000011 | -16.953125)   => (110.01111 | -1.53125)        
    3012 => 207,          -- (101111.000100 | -16.9375)     => (110.01111 | -1.53125)        
    3013 => 207,          -- (101111.000101 | -16.921875)   => (110.01111 | -1.53125)        
    3014 => 207,          -- (101111.000110 | -16.90625)    => (110.01111 | -1.53125)        
    3015 => 207,          -- (101111.000111 | -16.890625)   => (110.01111 | -1.53125)        
    3016 => 207,          -- (101111.001000 | -16.875)      => (110.01111 | -1.53125)        
    3017 => 207,          -- (101111.001001 | -16.859375)   => (110.01111 | -1.53125)        
    3018 => 207,          -- (101111.001010 | -16.84375)    => (110.01111 | -1.53125)        
    3019 => 207,          -- (101111.001011 | -16.828125)   => (110.01111 | -1.53125)        
    3020 => 207,          -- (101111.001100 | -16.8125)     => (110.01111 | -1.53125)        
    3021 => 207,          -- (101111.001101 | -16.796875)   => (110.01111 | -1.53125)        
    3022 => 207,          -- (101111.001110 | -16.78125)    => (110.01111 | -1.53125)        
    3023 => 207,          -- (101111.001111 | -16.765625)   => (110.01111 | -1.53125)        
    3024 => 207,          -- (101111.010000 | -16.75)       => (110.01111 | -1.53125)        
    3025 => 207,          -- (101111.010001 | -16.734375)   => (110.01111 | -1.53125)        
    3026 => 207,          -- (101111.010010 | -16.71875)    => (110.01111 | -1.53125)        
    3027 => 207,          -- (101111.010011 | -16.703125)   => (110.01111 | -1.53125)        
    3028 => 207,          -- (101111.010100 | -16.6875)     => (110.01111 | -1.53125)        
    3029 => 207,          -- (101111.010101 | -16.671875)   => (110.01111 | -1.53125)        
    3030 => 207,          -- (101111.010110 | -16.65625)    => (110.01111 | -1.53125)        
    3031 => 207,          -- (101111.010111 | -16.640625)   => (110.01111 | -1.53125)        
    3032 => 207,          -- (101111.011000 | -16.625)      => (110.01111 | -1.53125)        
    3033 => 207,          -- (101111.011001 | -16.609375)   => (110.01111 | -1.53125)        
    3034 => 207,          -- (101111.011010 | -16.59375)    => (110.01111 | -1.53125)        
    3035 => 207,          -- (101111.011011 | -16.578125)   => (110.01111 | -1.53125)        
    3036 => 207,          -- (101111.011100 | -16.5625)     => (110.01111 | -1.53125)        
    3037 => 207,          -- (101111.011101 | -16.546875)   => (110.01111 | -1.53125)        
    3038 => 207,          -- (101111.011110 | -16.53125)    => (110.01111 | -1.53125)        
    3039 => 207,          -- (101111.011111 | -16.515625)   => (110.01111 | -1.53125)        
    3040 => 207,          -- (101111.100000 | -16.5)        => (110.01111 | -1.53125)        
    3041 => 207,          -- (101111.100001 | -16.484375)   => (110.01111 | -1.53125)        
    3042 => 207,          -- (101111.100010 | -16.46875)    => (110.01111 | -1.53125)        
    3043 => 207,          -- (101111.100011 | -16.453125)   => (110.01111 | -1.53125)        
    3044 => 207,          -- (101111.100100 | -16.4375)     => (110.01111 | -1.53125)        
    3045 => 207,          -- (101111.100101 | -16.421875)   => (110.01111 | -1.53125)        
    3046 => 207,          -- (101111.100110 | -16.40625)    => (110.01111 | -1.53125)        
    3047 => 207,          -- (101111.100111 | -16.390625)   => (110.01111 | -1.53125)        
    3048 => 207,          -- (101111.101000 | -16.375)      => (110.01111 | -1.53125)        
    3049 => 207,          -- (101111.101001 | -16.359375)   => (110.01111 | -1.53125)        
    3050 => 207,          -- (101111.101010 | -16.34375)    => (110.01111 | -1.53125)        
    3051 => 207,          -- (101111.101011 | -16.328125)   => (110.01111 | -1.53125)        
    3052 => 207,          -- (101111.101100 | -16.3125)     => (110.01111 | -1.53125)        
    3053 => 207,          -- (101111.101101 | -16.296875)   => (110.01111 | -1.53125)        
    3054 => 207,          -- (101111.101110 | -16.28125)    => (110.01111 | -1.53125)        
    3055 => 207,          -- (101111.101111 | -16.265625)   => (110.01111 | -1.53125)        
    3056 => 207,          -- (101111.110000 | -16.25)       => (110.01111 | -1.53125)        
    3057 => 207,          -- (101111.110001 | -16.234375)   => (110.01111 | -1.53125)        
    3058 => 207,          -- (101111.110010 | -16.21875)    => (110.01111 | -1.53125)        
    3059 => 207,          -- (101111.110011 | -16.203125)   => (110.01111 | -1.53125)        
    3060 => 207,          -- (101111.110100 | -16.1875)     => (110.01111 | -1.53125)        
    3061 => 207,          -- (101111.110101 | -16.171875)   => (110.01111 | -1.53125)        
    3062 => 207,          -- (101111.110110 | -16.15625)    => (110.01111 | -1.53125)        
    3063 => 207,          -- (101111.110111 | -16.140625)   => (110.01111 | -1.53125)        
    3064 => 207,          -- (101111.111000 | -16.125)      => (110.01111 | -1.53125)        
    3065 => 207,          -- (101111.111001 | -16.109375)   => (110.01111 | -1.53125)        
    3066 => 207,          -- (101111.111010 | -16.09375)    => (110.01111 | -1.53125)        
    3067 => 207,          -- (101111.111011 | -16.078125)   => (110.01111 | -1.53125)        
    3068 => 207,          -- (101111.111100 | -16.0625)     => (110.01111 | -1.53125)        
    3069 => 207,          -- (101111.111101 | -16.046875)   => (110.01111 | -1.53125)        
    3070 => 207,          -- (101111.111110 | -16.03125)    => (110.01111 | -1.53125)        
    3071 => 207,          -- (101111.111111 | -16.015625)   => (110.01111 | -1.53125)        
    3072 => 207,          -- (110000.000000 | -16.0)        => (110.01111 | -1.53125)        
    3073 => 207,          -- (110000.000001 | -15.984375)   => (110.01111 | -1.53125)        
    3074 => 207,          -- (110000.000010 | -15.96875)    => (110.01111 | -1.53125)        
    3075 => 207,          -- (110000.000011 | -15.953125)   => (110.01111 | -1.53125)        
    3076 => 207,          -- (110000.000100 | -15.9375)     => (110.01111 | -1.53125)        
    3077 => 207,          -- (110000.000101 | -15.921875)   => (110.01111 | -1.53125)        
    3078 => 207,          -- (110000.000110 | -15.90625)    => (110.01111 | -1.53125)        
    3079 => 207,          -- (110000.000111 | -15.890625)   => (110.01111 | -1.53125)        
    3080 => 207,          -- (110000.001000 | -15.875)      => (110.01111 | -1.53125)        
    3081 => 207,          -- (110000.001001 | -15.859375)   => (110.01111 | -1.53125)        
    3082 => 207,          -- (110000.001010 | -15.84375)    => (110.01111 | -1.53125)        
    3083 => 207,          -- (110000.001011 | -15.828125)   => (110.01111 | -1.53125)        
    3084 => 207,          -- (110000.001100 | -15.8125)     => (110.01111 | -1.53125)        
    3085 => 207,          -- (110000.001101 | -15.796875)   => (110.01111 | -1.53125)        
    3086 => 207,          -- (110000.001110 | -15.78125)    => (110.01111 | -1.53125)        
    3087 => 207,          -- (110000.001111 | -15.765625)   => (110.01111 | -1.53125)        
    3088 => 207,          -- (110000.010000 | -15.75)       => (110.01111 | -1.53125)        
    3089 => 207,          -- (110000.010001 | -15.734375)   => (110.01111 | -1.53125)        
    3090 => 207,          -- (110000.010010 | -15.71875)    => (110.01111 | -1.53125)        
    3091 => 207,          -- (110000.010011 | -15.703125)   => (110.01111 | -1.53125)        
    3092 => 207,          -- (110000.010100 | -15.6875)     => (110.01111 | -1.53125)        
    3093 => 207,          -- (110000.010101 | -15.671875)   => (110.01111 | -1.53125)        
    3094 => 207,          -- (110000.010110 | -15.65625)    => (110.01111 | -1.53125)        
    3095 => 207,          -- (110000.010111 | -15.640625)   => (110.01111 | -1.53125)        
    3096 => 207,          -- (110000.011000 | -15.625)      => (110.01111 | -1.53125)        
    3097 => 207,          -- (110000.011001 | -15.609375)   => (110.01111 | -1.53125)        
    3098 => 207,          -- (110000.011010 | -15.59375)    => (110.01111 | -1.53125)        
    3099 => 207,          -- (110000.011011 | -15.578125)   => (110.01111 | -1.53125)        
    3100 => 207,          -- (110000.011100 | -15.5625)     => (110.01111 | -1.53125)        
    3101 => 207,          -- (110000.011101 | -15.546875)   => (110.01111 | -1.53125)        
    3102 => 207,          -- (110000.011110 | -15.53125)    => (110.01111 | -1.53125)        
    3103 => 207,          -- (110000.011111 | -15.515625)   => (110.01111 | -1.53125)        
    3104 => 207,          -- (110000.100000 | -15.5)        => (110.01111 | -1.53125)        
    3105 => 207,          -- (110000.100001 | -15.484375)   => (110.01111 | -1.53125)        
    3106 => 207,          -- (110000.100010 | -15.46875)    => (110.01111 | -1.53125)        
    3107 => 207,          -- (110000.100011 | -15.453125)   => (110.01111 | -1.53125)        
    3108 => 207,          -- (110000.100100 | -15.4375)     => (110.01111 | -1.53125)        
    3109 => 207,          -- (110000.100101 | -15.421875)   => (110.01111 | -1.53125)        
    3110 => 207,          -- (110000.100110 | -15.40625)    => (110.01111 | -1.53125)        
    3111 => 207,          -- (110000.100111 | -15.390625)   => (110.01111 | -1.53125)        
    3112 => 207,          -- (110000.101000 | -15.375)      => (110.01111 | -1.53125)        
    3113 => 207,          -- (110000.101001 | -15.359375)   => (110.01111 | -1.53125)        
    3114 => 207,          -- (110000.101010 | -15.34375)    => (110.01111 | -1.53125)        
    3115 => 207,          -- (110000.101011 | -15.328125)   => (110.01111 | -1.53125)        
    3116 => 207,          -- (110000.101100 | -15.3125)     => (110.01111 | -1.53125)        
    3117 => 207,          -- (110000.101101 | -15.296875)   => (110.01111 | -1.53125)        
    3118 => 207,          -- (110000.101110 | -15.28125)    => (110.01111 | -1.53125)        
    3119 => 207,          -- (110000.101111 | -15.265625)   => (110.01111 | -1.53125)        
    3120 => 207,          -- (110000.110000 | -15.25)       => (110.01111 | -1.53125)        
    3121 => 207,          -- (110000.110001 | -15.234375)   => (110.01111 | -1.53125)        
    3122 => 207,          -- (110000.110010 | -15.21875)    => (110.01111 | -1.53125)        
    3123 => 207,          -- (110000.110011 | -15.203125)   => (110.01111 | -1.53125)        
    3124 => 207,          -- (110000.110100 | -15.1875)     => (110.01111 | -1.53125)        
    3125 => 207,          -- (110000.110101 | -15.171875)   => (110.01111 | -1.53125)        
    3126 => 207,          -- (110000.110110 | -15.15625)    => (110.01111 | -1.53125)        
    3127 => 207,          -- (110000.110111 | -15.140625)   => (110.01111 | -1.53125)        
    3128 => 207,          -- (110000.111000 | -15.125)      => (110.01111 | -1.53125)        
    3129 => 207,          -- (110000.111001 | -15.109375)   => (110.01111 | -1.53125)        
    3130 => 207,          -- (110000.111010 | -15.09375)    => (110.01111 | -1.53125)        
    3131 => 207,          -- (110000.111011 | -15.078125)   => (110.01111 | -1.53125)        
    3132 => 207,          -- (110000.111100 | -15.0625)     => (110.01111 | -1.53125)        
    3133 => 207,          -- (110000.111101 | -15.046875)   => (110.01111 | -1.53125)        
    3134 => 207,          -- (110000.111110 | -15.03125)    => (110.01111 | -1.53125)        
    3135 => 207,          -- (110000.111111 | -15.015625)   => (110.01111 | -1.53125)        
    3136 => 207,          -- (110001.000000 | -15.0)        => (110.01111 | -1.53125)        
    3137 => 207,          -- (110001.000001 | -14.984375)   => (110.01111 | -1.53125)        
    3138 => 207,          -- (110001.000010 | -14.96875)    => (110.01111 | -1.53125)        
    3139 => 207,          -- (110001.000011 | -14.953125)   => (110.01111 | -1.53125)        
    3140 => 207,          -- (110001.000100 | -14.9375)     => (110.01111 | -1.53125)        
    3141 => 207,          -- (110001.000101 | -14.921875)   => (110.01111 | -1.53125)        
    3142 => 207,          -- (110001.000110 | -14.90625)    => (110.01111 | -1.53125)        
    3143 => 207,          -- (110001.000111 | -14.890625)   => (110.01111 | -1.53125)        
    3144 => 207,          -- (110001.001000 | -14.875)      => (110.01111 | -1.53125)        
    3145 => 207,          -- (110001.001001 | -14.859375)   => (110.01111 | -1.53125)        
    3146 => 207,          -- (110001.001010 | -14.84375)    => (110.01111 | -1.53125)        
    3147 => 207,          -- (110001.001011 | -14.828125)   => (110.01111 | -1.53125)        
    3148 => 207,          -- (110001.001100 | -14.8125)     => (110.01111 | -1.53125)        
    3149 => 207,          -- (110001.001101 | -14.796875)   => (110.01111 | -1.53125)        
    3150 => 207,          -- (110001.001110 | -14.78125)    => (110.01111 | -1.53125)        
    3151 => 207,          -- (110001.001111 | -14.765625)   => (110.01111 | -1.53125)        
    3152 => 207,          -- (110001.010000 | -14.75)       => (110.01111 | -1.53125)        
    3153 => 207,          -- (110001.010001 | -14.734375)   => (110.01111 | -1.53125)        
    3154 => 207,          -- (110001.010010 | -14.71875)    => (110.01111 | -1.53125)        
    3155 => 207,          -- (110001.010011 | -14.703125)   => (110.01111 | -1.53125)        
    3156 => 207,          -- (110001.010100 | -14.6875)     => (110.01111 | -1.53125)        
    3157 => 207,          -- (110001.010101 | -14.671875)   => (110.01111 | -1.53125)        
    3158 => 207,          -- (110001.010110 | -14.65625)    => (110.01111 | -1.53125)        
    3159 => 207,          -- (110001.010111 | -14.640625)   => (110.01111 | -1.53125)        
    3160 => 207,          -- (110001.011000 | -14.625)      => (110.01111 | -1.53125)        
    3161 => 207,          -- (110001.011001 | -14.609375)   => (110.01111 | -1.53125)        
    3162 => 207,          -- (110001.011010 | -14.59375)    => (110.01111 | -1.53125)        
    3163 => 207,          -- (110001.011011 | -14.578125)   => (110.01111 | -1.53125)        
    3164 => 207,          -- (110001.011100 | -14.5625)     => (110.01111 | -1.53125)        
    3165 => 207,          -- (110001.011101 | -14.546875)   => (110.01111 | -1.53125)        
    3166 => 207,          -- (110001.011110 | -14.53125)    => (110.01111 | -1.53125)        
    3167 => 207,          -- (110001.011111 | -14.515625)   => (110.01111 | -1.53125)        
    3168 => 207,          -- (110001.100000 | -14.5)        => (110.01111 | -1.53125)        
    3169 => 207,          -- (110001.100001 | -14.484375)   => (110.01111 | -1.53125)        
    3170 => 207,          -- (110001.100010 | -14.46875)    => (110.01111 | -1.53125)        
    3171 => 207,          -- (110001.100011 | -14.453125)   => (110.01111 | -1.53125)        
    3172 => 207,          -- (110001.100100 | -14.4375)     => (110.01111 | -1.53125)        
    3173 => 207,          -- (110001.100101 | -14.421875)   => (110.01111 | -1.53125)        
    3174 => 207,          -- (110001.100110 | -14.40625)    => (110.01111 | -1.53125)        
    3175 => 207,          -- (110001.100111 | -14.390625)   => (110.01111 | -1.53125)        
    3176 => 207,          -- (110001.101000 | -14.375)      => (110.01111 | -1.53125)        
    3177 => 207,          -- (110001.101001 | -14.359375)   => (110.01111 | -1.53125)        
    3178 => 207,          -- (110001.101010 | -14.34375)    => (110.01111 | -1.53125)        
    3179 => 207,          -- (110001.101011 | -14.328125)   => (110.01111 | -1.53125)        
    3180 => 207,          -- (110001.101100 | -14.3125)     => (110.01111 | -1.53125)        
    3181 => 207,          -- (110001.101101 | -14.296875)   => (110.01111 | -1.53125)        
    3182 => 207,          -- (110001.101110 | -14.28125)    => (110.01111 | -1.53125)        
    3183 => 207,          -- (110001.101111 | -14.265625)   => (110.01111 | -1.53125)        
    3184 => 207,          -- (110001.110000 | -14.25)       => (110.01111 | -1.53125)        
    3185 => 207,          -- (110001.110001 | -14.234375)   => (110.01111 | -1.53125)        
    3186 => 207,          -- (110001.110010 | -14.21875)    => (110.01111 | -1.53125)        
    3187 => 207,          -- (110001.110011 | -14.203125)   => (110.01111 | -1.53125)        
    3188 => 207,          -- (110001.110100 | -14.1875)     => (110.01111 | -1.53125)        
    3189 => 207,          -- (110001.110101 | -14.171875)   => (110.01111 | -1.53125)        
    3190 => 207,          -- (110001.110110 | -14.15625)    => (110.01111 | -1.53125)        
    3191 => 207,          -- (110001.110111 | -14.140625)   => (110.01111 | -1.53125)        
    3192 => 207,          -- (110001.111000 | -14.125)      => (110.01111 | -1.53125)        
    3193 => 207,          -- (110001.111001 | -14.109375)   => (110.01111 | -1.53125)        
    3194 => 208,          -- (110001.111010 | -14.09375)    => (110.10000 | -1.5)            
    3195 => 208,          -- (110001.111011 | -14.078125)   => (110.10000 | -1.5)            
    3196 => 208,          -- (110001.111100 | -14.0625)     => (110.10000 | -1.5)            
    3197 => 208,          -- (110001.111101 | -14.046875)   => (110.10000 | -1.5)            
    3198 => 208,          -- (110001.111110 | -14.03125)    => (110.10000 | -1.5)            
    3199 => 208,          -- (110001.111111 | -14.015625)   => (110.10000 | -1.5)            
    3200 => 208,          -- (110010.000000 | -14.0)        => (110.10000 | -1.5)            
    3201 => 208,          -- (110010.000001 | -13.984375)   => (110.10000 | -1.5)            
    3202 => 208,          -- (110010.000010 | -13.96875)    => (110.10000 | -1.5)            
    3203 => 208,          -- (110010.000011 | -13.953125)   => (110.10000 | -1.5)            
    3204 => 208,          -- (110010.000100 | -13.9375)     => (110.10000 | -1.5)            
    3205 => 208,          -- (110010.000101 | -13.921875)   => (110.10000 | -1.5)            
    3206 => 208,          -- (110010.000110 | -13.90625)    => (110.10000 | -1.5)            
    3207 => 208,          -- (110010.000111 | -13.890625)   => (110.10000 | -1.5)            
    3208 => 208,          -- (110010.001000 | -13.875)      => (110.10000 | -1.5)            
    3209 => 208,          -- (110010.001001 | -13.859375)   => (110.10000 | -1.5)            
    3210 => 208,          -- (110010.001010 | -13.84375)    => (110.10000 | -1.5)            
    3211 => 208,          -- (110010.001011 | -13.828125)   => (110.10000 | -1.5)            
    3212 => 208,          -- (110010.001100 | -13.8125)     => (110.10000 | -1.5)            
    3213 => 208,          -- (110010.001101 | -13.796875)   => (110.10000 | -1.5)            
    3214 => 208,          -- (110010.001110 | -13.78125)    => (110.10000 | -1.5)            
    3215 => 208,          -- (110010.001111 | -13.765625)   => (110.10000 | -1.5)            
    3216 => 208,          -- (110010.010000 | -13.75)       => (110.10000 | -1.5)            
    3217 => 208,          -- (110010.010001 | -13.734375)   => (110.10000 | -1.5)            
    3218 => 208,          -- (110010.010010 | -13.71875)    => (110.10000 | -1.5)            
    3219 => 208,          -- (110010.010011 | -13.703125)   => (110.10000 | -1.5)            
    3220 => 208,          -- (110010.010100 | -13.6875)     => (110.10000 | -1.5)            
    3221 => 208,          -- (110010.010101 | -13.671875)   => (110.10000 | -1.5)            
    3222 => 208,          -- (110010.010110 | -13.65625)    => (110.10000 | -1.5)            
    3223 => 208,          -- (110010.010111 | -13.640625)   => (110.10000 | -1.5)            
    3224 => 208,          -- (110010.011000 | -13.625)      => (110.10000 | -1.5)            
    3225 => 208,          -- (110010.011001 | -13.609375)   => (110.10000 | -1.5)            
    3226 => 208,          -- (110010.011010 | -13.59375)    => (110.10000 | -1.5)            
    3227 => 208,          -- (110010.011011 | -13.578125)   => (110.10000 | -1.5)            
    3228 => 208,          -- (110010.011100 | -13.5625)     => (110.10000 | -1.5)            
    3229 => 208,          -- (110010.011101 | -13.546875)   => (110.10000 | -1.5)            
    3230 => 208,          -- (110010.011110 | -13.53125)    => (110.10000 | -1.5)            
    3231 => 208,          -- (110010.011111 | -13.515625)   => (110.10000 | -1.5)            
    3232 => 208,          -- (110010.100000 | -13.5)        => (110.10000 | -1.5)            
    3233 => 208,          -- (110010.100001 | -13.484375)   => (110.10000 | -1.5)            
    3234 => 208,          -- (110010.100010 | -13.46875)    => (110.10000 | -1.5)            
    3235 => 208,          -- (110010.100011 | -13.453125)   => (110.10000 | -1.5)            
    3236 => 208,          -- (110010.100100 | -13.4375)     => (110.10000 | -1.5)            
    3237 => 208,          -- (110010.100101 | -13.421875)   => (110.10000 | -1.5)            
    3238 => 208,          -- (110010.100110 | -13.40625)    => (110.10000 | -1.5)            
    3239 => 208,          -- (110010.100111 | -13.390625)   => (110.10000 | -1.5)            
    3240 => 208,          -- (110010.101000 | -13.375)      => (110.10000 | -1.5)            
    3241 => 208,          -- (110010.101001 | -13.359375)   => (110.10000 | -1.5)            
    3242 => 208,          -- (110010.101010 | -13.34375)    => (110.10000 | -1.5)            
    3243 => 208,          -- (110010.101011 | -13.328125)   => (110.10000 | -1.5)            
    3244 => 208,          -- (110010.101100 | -13.3125)     => (110.10000 | -1.5)            
    3245 => 208,          -- (110010.101101 | -13.296875)   => (110.10000 | -1.5)            
    3246 => 208,          -- (110010.101110 | -13.28125)    => (110.10000 | -1.5)            
    3247 => 208,          -- (110010.101111 | -13.265625)   => (110.10000 | -1.5)            
    3248 => 208,          -- (110010.110000 | -13.25)       => (110.10000 | -1.5)            
    3249 => 208,          -- (110010.110001 | -13.234375)   => (110.10000 | -1.5)            
    3250 => 208,          -- (110010.110010 | -13.21875)    => (110.10000 | -1.5)            
    3251 => 208,          -- (110010.110011 | -13.203125)   => (110.10000 | -1.5)            
    3252 => 208,          -- (110010.110100 | -13.1875)     => (110.10000 | -1.5)            
    3253 => 208,          -- (110010.110101 | -13.171875)   => (110.10000 | -1.5)            
    3254 => 208,          -- (110010.110110 | -13.15625)    => (110.10000 | -1.5)            
    3255 => 208,          -- (110010.110111 | -13.140625)   => (110.10000 | -1.5)            
    3256 => 208,          -- (110010.111000 | -13.125)      => (110.10000 | -1.5)            
    3257 => 208,          -- (110010.111001 | -13.109375)   => (110.10000 | -1.5)            
    3258 => 208,          -- (110010.111010 | -13.09375)    => (110.10000 | -1.5)            
    3259 => 208,          -- (110010.111011 | -13.078125)   => (110.10000 | -1.5)            
    3260 => 208,          -- (110010.111100 | -13.0625)     => (110.10000 | -1.5)            
    3261 => 208,          -- (110010.111101 | -13.046875)   => (110.10000 | -1.5)            
    3262 => 208,          -- (110010.111110 | -13.03125)    => (110.10000 | -1.5)            
    3263 => 208,          -- (110010.111111 | -13.015625)   => (110.10000 | -1.5)            
    3264 => 208,          -- (110011.000000 | -13.0)        => (110.10000 | -1.5)            
    3265 => 208,          -- (110011.000001 | -12.984375)   => (110.10000 | -1.5)            
    3266 => 208,          -- (110011.000010 | -12.96875)    => (110.10000 | -1.5)            
    3267 => 208,          -- (110011.000011 | -12.953125)   => (110.10000 | -1.5)            
    3268 => 208,          -- (110011.000100 | -12.9375)     => (110.10000 | -1.5)            
    3269 => 208,          -- (110011.000101 | -12.921875)   => (110.10000 | -1.5)            
    3270 => 208,          -- (110011.000110 | -12.90625)    => (110.10000 | -1.5)            
    3271 => 208,          -- (110011.000111 | -12.890625)   => (110.10000 | -1.5)            
    3272 => 208,          -- (110011.001000 | -12.875)      => (110.10000 | -1.5)            
    3273 => 208,          -- (110011.001001 | -12.859375)   => (110.10000 | -1.5)            
    3274 => 208,          -- (110011.001010 | -12.84375)    => (110.10000 | -1.5)            
    3275 => 208,          -- (110011.001011 | -12.828125)   => (110.10000 | -1.5)            
    3276 => 208,          -- (110011.001100 | -12.8125)     => (110.10000 | -1.5)            
    3277 => 208,          -- (110011.001101 | -12.796875)   => (110.10000 | -1.5)            
    3278 => 208,          -- (110011.001110 | -12.78125)    => (110.10000 | -1.5)            
    3279 => 208,          -- (110011.001111 | -12.765625)   => (110.10000 | -1.5)            
    3280 => 208,          -- (110011.010000 | -12.75)       => (110.10000 | -1.5)            
    3281 => 208,          -- (110011.010001 | -12.734375)   => (110.10000 | -1.5)            
    3282 => 208,          -- (110011.010010 | -12.71875)    => (110.10000 | -1.5)            
    3283 => 208,          -- (110011.010011 | -12.703125)   => (110.10000 | -1.5)            
    3284 => 208,          -- (110011.010100 | -12.6875)     => (110.10000 | -1.5)            
    3285 => 208,          -- (110011.010101 | -12.671875)   => (110.10000 | -1.5)            
    3286 => 208,          -- (110011.010110 | -12.65625)    => (110.10000 | -1.5)            
    3287 => 208,          -- (110011.010111 | -12.640625)   => (110.10000 | -1.5)            
    3288 => 208,          -- (110011.011000 | -12.625)      => (110.10000 | -1.5)            
    3289 => 208,          -- (110011.011001 | -12.609375)   => (110.10000 | -1.5)            
    3290 => 208,          -- (110011.011010 | -12.59375)    => (110.10000 | -1.5)            
    3291 => 208,          -- (110011.011011 | -12.578125)   => (110.10000 | -1.5)            
    3292 => 208,          -- (110011.011100 | -12.5625)     => (110.10000 | -1.5)            
    3293 => 208,          -- (110011.011101 | -12.546875)   => (110.10000 | -1.5)            
    3294 => 208,          -- (110011.011110 | -12.53125)    => (110.10000 | -1.5)            
    3295 => 208,          -- (110011.011111 | -12.515625)   => (110.10000 | -1.5)            
    3296 => 208,          -- (110011.100000 | -12.5)        => (110.10000 | -1.5)            
    3297 => 208,          -- (110011.100001 | -12.484375)   => (110.10000 | -1.5)            
    3298 => 208,          -- (110011.100010 | -12.46875)    => (110.10000 | -1.5)            
    3299 => 208,          -- (110011.100011 | -12.453125)   => (110.10000 | -1.5)            
    3300 => 208,          -- (110011.100100 | -12.4375)     => (110.10000 | -1.5)            
    3301 => 208,          -- (110011.100101 | -12.421875)   => (110.10000 | -1.5)            
    3302 => 208,          -- (110011.100110 | -12.40625)    => (110.10000 | -1.5)            
    3303 => 208,          -- (110011.100111 | -12.390625)   => (110.10000 | -1.5)            
    3304 => 208,          -- (110011.101000 | -12.375)      => (110.10000 | -1.5)            
    3305 => 208,          -- (110011.101001 | -12.359375)   => (110.10000 | -1.5)            
    3306 => 208,          -- (110011.101010 | -12.34375)    => (110.10000 | -1.5)            
    3307 => 208,          -- (110011.101011 | -12.328125)   => (110.10000 | -1.5)            
    3308 => 208,          -- (110011.101100 | -12.3125)     => (110.10000 | -1.5)            
    3309 => 208,          -- (110011.101101 | -12.296875)   => (110.10000 | -1.5)            
    3310 => 208,          -- (110011.101110 | -12.28125)    => (110.10000 | -1.5)            
    3311 => 208,          -- (110011.101111 | -12.265625)   => (110.10000 | -1.5)            
    3312 => 208,          -- (110011.110000 | -12.25)       => (110.10000 | -1.5)            
    3313 => 208,          -- (110011.110001 | -12.234375)   => (110.10000 | -1.5)            
    3314 => 208,          -- (110011.110010 | -12.21875)    => (110.10000 | -1.5)            
    3315 => 208,          -- (110011.110011 | -12.203125)   => (110.10000 | -1.5)            
    3316 => 208,          -- (110011.110100 | -12.1875)     => (110.10000 | -1.5)            
    3317 => 208,          -- (110011.110101 | -12.171875)   => (110.10000 | -1.5)            
    3318 => 208,          -- (110011.110110 | -12.15625)    => (110.10000 | -1.5)            
    3319 => 208,          -- (110011.110111 | -12.140625)   => (110.10000 | -1.5)            
    3320 => 208,          -- (110011.111000 | -12.125)      => (110.10000 | -1.5)            
    3321 => 208,          -- (110011.111001 | -12.109375)   => (110.10000 | -1.5)            
    3322 => 208,          -- (110011.111010 | -12.09375)    => (110.10000 | -1.5)            
    3323 => 208,          -- (110011.111011 | -12.078125)   => (110.10000 | -1.5)            
    3324 => 208,          -- (110011.111100 | -12.0625)     => (110.10000 | -1.5)            
    3325 => 208,          -- (110011.111101 | -12.046875)   => (110.10000 | -1.5)            
    3326 => 208,          -- (110011.111110 | -12.03125)    => (110.10000 | -1.5)            
    3327 => 208,          -- (110011.111111 | -12.015625)   => (110.10000 | -1.5)            
    3328 => 208,          -- (110100.000000 | -12.0)        => (110.10000 | -1.5)            
    3329 => 208,          -- (110100.000001 | -11.984375)   => (110.10000 | -1.5)            
    3330 => 208,          -- (110100.000010 | -11.96875)    => (110.10000 | -1.5)            
    3331 => 208,          -- (110100.000011 | -11.953125)   => (110.10000 | -1.5)            
    3332 => 208,          -- (110100.000100 | -11.9375)     => (110.10000 | -1.5)            
    3333 => 208,          -- (110100.000101 | -11.921875)   => (110.10000 | -1.5)            
    3334 => 208,          -- (110100.000110 | -11.90625)    => (110.10000 | -1.5)            
    3335 => 208,          -- (110100.000111 | -11.890625)   => (110.10000 | -1.5)            
    3336 => 208,          -- (110100.001000 | -11.875)      => (110.10000 | -1.5)            
    3337 => 208,          -- (110100.001001 | -11.859375)   => (110.10000 | -1.5)            
    3338 => 208,          -- (110100.001010 | -11.84375)    => (110.10000 | -1.5)            
    3339 => 208,          -- (110100.001011 | -11.828125)   => (110.10000 | -1.5)            
    3340 => 208,          -- (110100.001100 | -11.8125)     => (110.10000 | -1.5)            
    3341 => 208,          -- (110100.001101 | -11.796875)   => (110.10000 | -1.5)            
    3342 => 208,          -- (110100.001110 | -11.78125)    => (110.10000 | -1.5)            
    3343 => 208,          -- (110100.001111 | -11.765625)   => (110.10000 | -1.5)            
    3344 => 208,          -- (110100.010000 | -11.75)       => (110.10000 | -1.5)            
    3345 => 208,          -- (110100.010001 | -11.734375)   => (110.10000 | -1.5)            
    3346 => 208,          -- (110100.010010 | -11.71875)    => (110.10000 | -1.5)            
    3347 => 208,          -- (110100.010011 | -11.703125)   => (110.10000 | -1.5)            
    3348 => 208,          -- (110100.010100 | -11.6875)     => (110.10000 | -1.5)            
    3349 => 208,          -- (110100.010101 | -11.671875)   => (110.10000 | -1.5)            
    3350 => 208,          -- (110100.010110 | -11.65625)    => (110.10000 | -1.5)            
    3351 => 208,          -- (110100.010111 | -11.640625)   => (110.10000 | -1.5)            
    3352 => 208,          -- (110100.011000 | -11.625)      => (110.10000 | -1.5)            
    3353 => 208,          -- (110100.011001 | -11.609375)   => (110.10000 | -1.5)            
    3354 => 208,          -- (110100.011010 | -11.59375)    => (110.10000 | -1.5)            
    3355 => 208,          -- (110100.011011 | -11.578125)   => (110.10000 | -1.5)            
    3356 => 208,          -- (110100.011100 | -11.5625)     => (110.10000 | -1.5)            
    3357 => 208,          -- (110100.011101 | -11.546875)   => (110.10000 | -1.5)            
    3358 => 208,          -- (110100.011110 | -11.53125)    => (110.10000 | -1.5)            
    3359 => 208,          -- (110100.011111 | -11.515625)   => (110.10000 | -1.5)            
    3360 => 208,          -- (110100.100000 | -11.5)        => (110.10000 | -1.5)            
    3361 => 208,          -- (110100.100001 | -11.484375)   => (110.10000 | -1.5)            
    3362 => 208,          -- (110100.100010 | -11.46875)    => (110.10000 | -1.5)            
    3363 => 208,          -- (110100.100011 | -11.453125)   => (110.10000 | -1.5)            
    3364 => 208,          -- (110100.100100 | -11.4375)     => (110.10000 | -1.5)            
    3365 => 208,          -- (110100.100101 | -11.421875)   => (110.10000 | -1.5)            
    3366 => 208,          -- (110100.100110 | -11.40625)    => (110.10000 | -1.5)            
    3367 => 208,          -- (110100.100111 | -11.390625)   => (110.10000 | -1.5)            
    3368 => 208,          -- (110100.101000 | -11.375)      => (110.10000 | -1.5)            
    3369 => 208,          -- (110100.101001 | -11.359375)   => (110.10000 | -1.5)            
    3370 => 208,          -- (110100.101010 | -11.34375)    => (110.10000 | -1.5)            
    3371 => 208,          -- (110100.101011 | -11.328125)   => (110.10000 | -1.5)            
    3372 => 208,          -- (110100.101100 | -11.3125)     => (110.10000 | -1.5)            
    3373 => 208,          -- (110100.101101 | -11.296875)   => (110.10000 | -1.5)            
    3374 => 208,          -- (110100.101110 | -11.28125)    => (110.10000 | -1.5)            
    3375 => 208,          -- (110100.101111 | -11.265625)   => (110.10000 | -1.5)            
    3376 => 208,          -- (110100.110000 | -11.25)       => (110.10000 | -1.5)            
    3377 => 208,          -- (110100.110001 | -11.234375)   => (110.10000 | -1.5)            
    3378 => 208,          -- (110100.110010 | -11.21875)    => (110.10000 | -1.5)            
    3379 => 208,          -- (110100.110011 | -11.203125)   => (110.10000 | -1.5)            
    3380 => 208,          -- (110100.110100 | -11.1875)     => (110.10000 | -1.5)            
    3381 => 208,          -- (110100.110101 | -11.171875)   => (110.10000 | -1.5)            
    3382 => 208,          -- (110100.110110 | -11.15625)    => (110.10000 | -1.5)            
    3383 => 208,          -- (110100.110111 | -11.140625)   => (110.10000 | -1.5)            
    3384 => 208,          -- (110100.111000 | -11.125)      => (110.10000 | -1.5)            
    3385 => 208,          -- (110100.111001 | -11.109375)   => (110.10000 | -1.5)            
    3386 => 208,          -- (110100.111010 | -11.09375)    => (110.10000 | -1.5)            
    3387 => 208,          -- (110100.111011 | -11.078125)   => (110.10000 | -1.5)            
    3388 => 208,          -- (110100.111100 | -11.0625)     => (110.10000 | -1.5)            
    3389 => 208,          -- (110100.111101 | -11.046875)   => (110.10000 | -1.5)            
    3390 => 208,          -- (110100.111110 | -11.03125)    => (110.10000 | -1.5)            
    3391 => 208,          -- (110100.111111 | -11.015625)   => (110.10000 | -1.5)            
    3392 => 208,          -- (110101.000000 | -11.0)        => (110.10000 | -1.5)            
    3393 => 208,          -- (110101.000001 | -10.984375)   => (110.10000 | -1.5)            
    3394 => 208,          -- (110101.000010 | -10.96875)    => (110.10000 | -1.5)            
    3395 => 208,          -- (110101.000011 | -10.953125)   => (110.10000 | -1.5)            
    3396 => 208,          -- (110101.000100 | -10.9375)     => (110.10000 | -1.5)            
    3397 => 208,          -- (110101.000101 | -10.921875)   => (110.10000 | -1.5)            
    3398 => 208,          -- (110101.000110 | -10.90625)    => (110.10000 | -1.5)            
    3399 => 208,          -- (110101.000111 | -10.890625)   => (110.10000 | -1.5)            
    3400 => 208,          -- (110101.001000 | -10.875)      => (110.10000 | -1.5)            
    3401 => 208,          -- (110101.001001 | -10.859375)   => (110.10000 | -1.5)            
    3402 => 208,          -- (110101.001010 | -10.84375)    => (110.10000 | -1.5)            
    3403 => 208,          -- (110101.001011 | -10.828125)   => (110.10000 | -1.5)            
    3404 => 208,          -- (110101.001100 | -10.8125)     => (110.10000 | -1.5)            
    3405 => 208,          -- (110101.001101 | -10.796875)   => (110.10000 | -1.5)            
    3406 => 208,          -- (110101.001110 | -10.78125)    => (110.10000 | -1.5)            
    3407 => 208,          -- (110101.001111 | -10.765625)   => (110.10000 | -1.5)            
    3408 => 208,          -- (110101.010000 | -10.75)       => (110.10000 | -1.5)            
    3409 => 208,          -- (110101.010001 | -10.734375)   => (110.10000 | -1.5)            
    3410 => 208,          -- (110101.010010 | -10.71875)    => (110.10000 | -1.5)            
    3411 => 208,          -- (110101.010011 | -10.703125)   => (110.10000 | -1.5)            
    3412 => 208,          -- (110101.010100 | -10.6875)     => (110.10000 | -1.5)            
    3413 => 208,          -- (110101.010101 | -10.671875)   => (110.10000 | -1.5)            
    3414 => 208,          -- (110101.010110 | -10.65625)    => (110.10000 | -1.5)            
    3415 => 208,          -- (110101.010111 | -10.640625)   => (110.10000 | -1.5)            
    3416 => 208,          -- (110101.011000 | -10.625)      => (110.10000 | -1.5)            
    3417 => 208,          -- (110101.011001 | -10.609375)   => (110.10000 | -1.5)            
    3418 => 208,          -- (110101.011010 | -10.59375)    => (110.10000 | -1.5)            
    3419 => 208,          -- (110101.011011 | -10.578125)   => (110.10000 | -1.5)            
    3420 => 208,          -- (110101.011100 | -10.5625)     => (110.10000 | -1.5)            
    3421 => 208,          -- (110101.011101 | -10.546875)   => (110.10000 | -1.5)            
    3422 => 208,          -- (110101.011110 | -10.53125)    => (110.10000 | -1.5)            
    3423 => 208,          -- (110101.011111 | -10.515625)   => (110.10000 | -1.5)            
    3424 => 208,          -- (110101.100000 | -10.5)        => (110.10000 | -1.5)            
    3425 => 208,          -- (110101.100001 | -10.484375)   => (110.10000 | -1.5)            
    3426 => 208,          -- (110101.100010 | -10.46875)    => (110.10000 | -1.5)            
    3427 => 208,          -- (110101.100011 | -10.453125)   => (110.10000 | -1.5)            
    3428 => 208,          -- (110101.100100 | -10.4375)     => (110.10000 | -1.5)            
    3429 => 208,          -- (110101.100101 | -10.421875)   => (110.10000 | -1.5)            
    3430 => 208,          -- (110101.100110 | -10.40625)    => (110.10000 | -1.5)            
    3431 => 208,          -- (110101.100111 | -10.390625)   => (110.10000 | -1.5)            
    3432 => 208,          -- (110101.101000 | -10.375)      => (110.10000 | -1.5)            
    3433 => 208,          -- (110101.101001 | -10.359375)   => (110.10000 | -1.5)            
    3434 => 208,          -- (110101.101010 | -10.34375)    => (110.10000 | -1.5)            
    3435 => 208,          -- (110101.101011 | -10.328125)   => (110.10000 | -1.5)            
    3436 => 208,          -- (110101.101100 | -10.3125)     => (110.10000 | -1.5)            
    3437 => 208,          -- (110101.101101 | -10.296875)   => (110.10000 | -1.5)            
    3438 => 208,          -- (110101.101110 | -10.28125)    => (110.10000 | -1.5)            
    3439 => 208,          -- (110101.101111 | -10.265625)   => (110.10000 | -1.5)            
    3440 => 208,          -- (110101.110000 | -10.25)       => (110.10000 | -1.5)            
    3441 => 208,          -- (110101.110001 | -10.234375)   => (110.10000 | -1.5)            
    3442 => 208,          -- (110101.110010 | -10.21875)    => (110.10000 | -1.5)            
    3443 => 208,          -- (110101.110011 | -10.203125)   => (110.10000 | -1.5)            
    3444 => 208,          -- (110101.110100 | -10.1875)     => (110.10000 | -1.5)            
    3445 => 208,          -- (110101.110101 | -10.171875)   => (110.10000 | -1.5)            
    3446 => 208,          -- (110101.110110 | -10.15625)    => (110.10000 | -1.5)            
    3447 => 208,          -- (110101.110111 | -10.140625)   => (110.10000 | -1.5)            
    3448 => 208,          -- (110101.111000 | -10.125)      => (110.10000 | -1.5)            
    3449 => 208,          -- (110101.111001 | -10.109375)   => (110.10000 | -1.5)            
    3450 => 208,          -- (110101.111010 | -10.09375)    => (110.10000 | -1.5)            
    3451 => 208,          -- (110101.111011 | -10.078125)   => (110.10000 | -1.5)            
    3452 => 208,          -- (110101.111100 | -10.0625)     => (110.10000 | -1.5)            
    3453 => 208,          -- (110101.111101 | -10.046875)   => (110.10000 | -1.5)            
    3454 => 208,          -- (110101.111110 | -10.03125)    => (110.10000 | -1.5)            
    3455 => 208,          -- (110101.111111 | -10.015625)   => (110.10000 | -1.5)            
    3456 => 208,          -- (110110.000000 | -10.0)        => (110.10000 | -1.5)            
    3457 => 208,          -- (110110.000001 | -9.984375)    => (110.10000 | -1.5)            
    3458 => 208,          -- (110110.000010 | -9.96875)     => (110.10000 | -1.5)            
    3459 => 208,          -- (110110.000011 | -9.953125)    => (110.10000 | -1.5)            
    3460 => 208,          -- (110110.000100 | -9.9375)      => (110.10000 | -1.5)            
    3461 => 208,          -- (110110.000101 | -9.921875)    => (110.10000 | -1.5)            
    3462 => 208,          -- (110110.000110 | -9.90625)     => (110.10000 | -1.5)            
    3463 => 208,          -- (110110.000111 | -9.890625)    => (110.10000 | -1.5)            
    3464 => 208,          -- (110110.001000 | -9.875)       => (110.10000 | -1.5)            
    3465 => 208,          -- (110110.001001 | -9.859375)    => (110.10000 | -1.5)            
    3466 => 208,          -- (110110.001010 | -9.84375)     => (110.10000 | -1.5)            
    3467 => 208,          -- (110110.001011 | -9.828125)    => (110.10000 | -1.5)            
    3468 => 208,          -- (110110.001100 | -9.8125)      => (110.10000 | -1.5)            
    3469 => 208,          -- (110110.001101 | -9.796875)    => (110.10000 | -1.5)            
    3470 => 208,          -- (110110.001110 | -9.78125)     => (110.10000 | -1.5)            
    3471 => 208,          -- (110110.001111 | -9.765625)    => (110.10000 | -1.5)            
    3472 => 209,          -- (110110.010000 | -9.75)        => (110.10001 | -1.46875)        
    3473 => 209,          -- (110110.010001 | -9.734375)    => (110.10001 | -1.46875)        
    3474 => 209,          -- (110110.010010 | -9.71875)     => (110.10001 | -1.46875)        
    3475 => 209,          -- (110110.010011 | -9.703125)    => (110.10001 | -1.46875)        
    3476 => 209,          -- (110110.010100 | -9.6875)      => (110.10001 | -1.46875)        
    3477 => 209,          -- (110110.010101 | -9.671875)    => (110.10001 | -1.46875)        
    3478 => 209,          -- (110110.010110 | -9.65625)     => (110.10001 | -1.46875)        
    3479 => 209,          -- (110110.010111 | -9.640625)    => (110.10001 | -1.46875)        
    3480 => 209,          -- (110110.011000 | -9.625)       => (110.10001 | -1.46875)        
    3481 => 209,          -- (110110.011001 | -9.609375)    => (110.10001 | -1.46875)        
    3482 => 209,          -- (110110.011010 | -9.59375)     => (110.10001 | -1.46875)        
    3483 => 209,          -- (110110.011011 | -9.578125)    => (110.10001 | -1.46875)        
    3484 => 209,          -- (110110.011100 | -9.5625)      => (110.10001 | -1.46875)        
    3485 => 209,          -- (110110.011101 | -9.546875)    => (110.10001 | -1.46875)        
    3486 => 209,          -- (110110.011110 | -9.53125)     => (110.10001 | -1.46875)        
    3487 => 209,          -- (110110.011111 | -9.515625)    => (110.10001 | -1.46875)        
    3488 => 209,          -- (110110.100000 | -9.5)         => (110.10001 | -1.46875)        
    3489 => 209,          -- (110110.100001 | -9.484375)    => (110.10001 | -1.46875)        
    3490 => 209,          -- (110110.100010 | -9.46875)     => (110.10001 | -1.46875)        
    3491 => 209,          -- (110110.100011 | -9.453125)    => (110.10001 | -1.46875)        
    3492 => 209,          -- (110110.100100 | -9.4375)      => (110.10001 | -1.46875)        
    3493 => 209,          -- (110110.100101 | -9.421875)    => (110.10001 | -1.46875)        
    3494 => 209,          -- (110110.100110 | -9.40625)     => (110.10001 | -1.46875)        
    3495 => 209,          -- (110110.100111 | -9.390625)    => (110.10001 | -1.46875)        
    3496 => 209,          -- (110110.101000 | -9.375)       => (110.10001 | -1.46875)        
    3497 => 209,          -- (110110.101001 | -9.359375)    => (110.10001 | -1.46875)        
    3498 => 209,          -- (110110.101010 | -9.34375)     => (110.10001 | -1.46875)        
    3499 => 209,          -- (110110.101011 | -9.328125)    => (110.10001 | -1.46875)        
    3500 => 209,          -- (110110.101100 | -9.3125)      => (110.10001 | -1.46875)        
    3501 => 209,          -- (110110.101101 | -9.296875)    => (110.10001 | -1.46875)        
    3502 => 209,          -- (110110.101110 | -9.28125)     => (110.10001 | -1.46875)        
    3503 => 209,          -- (110110.101111 | -9.265625)    => (110.10001 | -1.46875)        
    3504 => 209,          -- (110110.110000 | -9.25)        => (110.10001 | -1.46875)        
    3505 => 209,          -- (110110.110001 | -9.234375)    => (110.10001 | -1.46875)        
    3506 => 209,          -- (110110.110010 | -9.21875)     => (110.10001 | -1.46875)        
    3507 => 209,          -- (110110.110011 | -9.203125)    => (110.10001 | -1.46875)        
    3508 => 209,          -- (110110.110100 | -9.1875)      => (110.10001 | -1.46875)        
    3509 => 209,          -- (110110.110101 | -9.171875)    => (110.10001 | -1.46875)        
    3510 => 209,          -- (110110.110110 | -9.15625)     => (110.10001 | -1.46875)        
    3511 => 209,          -- (110110.110111 | -9.140625)    => (110.10001 | -1.46875)        
    3512 => 209,          -- (110110.111000 | -9.125)       => (110.10001 | -1.46875)        
    3513 => 209,          -- (110110.111001 | -9.109375)    => (110.10001 | -1.46875)        
    3514 => 209,          -- (110110.111010 | -9.09375)     => (110.10001 | -1.46875)        
    3515 => 209,          -- (110110.111011 | -9.078125)    => (110.10001 | -1.46875)        
    3516 => 209,          -- (110110.111100 | -9.0625)      => (110.10001 | -1.46875)        
    3517 => 209,          -- (110110.111101 | -9.046875)    => (110.10001 | -1.46875)        
    3518 => 209,          -- (110110.111110 | -9.03125)     => (110.10001 | -1.46875)        
    3519 => 209,          -- (110110.111111 | -9.015625)    => (110.10001 | -1.46875)        
    3520 => 209,          -- (110111.000000 | -9.0)         => (110.10001 | -1.46875)        
    3521 => 209,          -- (110111.000001 | -8.984375)    => (110.10001 | -1.46875)        
    3522 => 209,          -- (110111.000010 | -8.96875)     => (110.10001 | -1.46875)        
    3523 => 209,          -- (110111.000011 | -8.953125)    => (110.10001 | -1.46875)        
    3524 => 209,          -- (110111.000100 | -8.9375)      => (110.10001 | -1.46875)        
    3525 => 209,          -- (110111.000101 | -8.921875)    => (110.10001 | -1.46875)        
    3526 => 209,          -- (110111.000110 | -8.90625)     => (110.10001 | -1.46875)        
    3527 => 209,          -- (110111.000111 | -8.890625)    => (110.10001 | -1.46875)        
    3528 => 209,          -- (110111.001000 | -8.875)       => (110.10001 | -1.46875)        
    3529 => 209,          -- (110111.001001 | -8.859375)    => (110.10001 | -1.46875)        
    3530 => 209,          -- (110111.001010 | -8.84375)     => (110.10001 | -1.46875)        
    3531 => 209,          -- (110111.001011 | -8.828125)    => (110.10001 | -1.46875)        
    3532 => 209,          -- (110111.001100 | -8.8125)      => (110.10001 | -1.46875)        
    3533 => 209,          -- (110111.001101 | -8.796875)    => (110.10001 | -1.46875)        
    3534 => 209,          -- (110111.001110 | -8.78125)     => (110.10001 | -1.46875)        
    3535 => 209,          -- (110111.001111 | -8.765625)    => (110.10001 | -1.46875)        
    3536 => 209,          -- (110111.010000 | -8.75)        => (110.10001 | -1.46875)        
    3537 => 209,          -- (110111.010001 | -8.734375)    => (110.10001 | -1.46875)        
    3538 => 209,          -- (110111.010010 | -8.71875)     => (110.10001 | -1.46875)        
    3539 => 209,          -- (110111.010011 | -8.703125)    => (110.10001 | -1.46875)        
    3540 => 209,          -- (110111.010100 | -8.6875)      => (110.10001 | -1.46875)        
    3541 => 209,          -- (110111.010101 | -8.671875)    => (110.10001 | -1.46875)        
    3542 => 209,          -- (110111.010110 | -8.65625)     => (110.10001 | -1.46875)        
    3543 => 209,          -- (110111.010111 | -8.640625)    => (110.10001 | -1.46875)        
    3544 => 209,          -- (110111.011000 | -8.625)       => (110.10001 | -1.46875)        
    3545 => 209,          -- (110111.011001 | -8.609375)    => (110.10001 | -1.46875)        
    3546 => 209,          -- (110111.011010 | -8.59375)     => (110.10001 | -1.46875)        
    3547 => 209,          -- (110111.011011 | -8.578125)    => (110.10001 | -1.46875)        
    3548 => 209,          -- (110111.011100 | -8.5625)      => (110.10001 | -1.46875)        
    3549 => 209,          -- (110111.011101 | -8.546875)    => (110.10001 | -1.46875)        
    3550 => 209,          -- (110111.011110 | -8.53125)     => (110.10001 | -1.46875)        
    3551 => 209,          -- (110111.011111 | -8.515625)    => (110.10001 | -1.46875)        
    3552 => 209,          -- (110111.100000 | -8.5)         => (110.10001 | -1.46875)        
    3553 => 209,          -- (110111.100001 | -8.484375)    => (110.10001 | -1.46875)        
    3554 => 209,          -- (110111.100010 | -8.46875)     => (110.10001 | -1.46875)        
    3555 => 209,          -- (110111.100011 | -8.453125)    => (110.10001 | -1.46875)        
    3556 => 209,          -- (110111.100100 | -8.4375)      => (110.10001 | -1.46875)        
    3557 => 209,          -- (110111.100101 | -8.421875)    => (110.10001 | -1.46875)        
    3558 => 209,          -- (110111.100110 | -8.40625)     => (110.10001 | -1.46875)        
    3559 => 209,          -- (110111.100111 | -8.390625)    => (110.10001 | -1.46875)        
    3560 => 209,          -- (110111.101000 | -8.375)       => (110.10001 | -1.46875)        
    3561 => 209,          -- (110111.101001 | -8.359375)    => (110.10001 | -1.46875)        
    3562 => 209,          -- (110111.101010 | -8.34375)     => (110.10001 | -1.46875)        
    3563 => 209,          -- (110111.101011 | -8.328125)    => (110.10001 | -1.46875)        
    3564 => 209,          -- (110111.101100 | -8.3125)      => (110.10001 | -1.46875)        
    3565 => 209,          -- (110111.101101 | -8.296875)    => (110.10001 | -1.46875)        
    3566 => 209,          -- (110111.101110 | -8.28125)     => (110.10001 | -1.46875)        
    3567 => 209,          -- (110111.101111 | -8.265625)    => (110.10001 | -1.46875)        
    3568 => 209,          -- (110111.110000 | -8.25)        => (110.10001 | -1.46875)        
    3569 => 209,          -- (110111.110001 | -8.234375)    => (110.10001 | -1.46875)        
    3570 => 209,          -- (110111.110010 | -8.21875)     => (110.10001 | -1.46875)        
    3571 => 209,          -- (110111.110011 | -8.203125)    => (110.10001 | -1.46875)        
    3572 => 209,          -- (110111.110100 | -8.1875)      => (110.10001 | -1.46875)        
    3573 => 209,          -- (110111.110101 | -8.171875)    => (110.10001 | -1.46875)        
    3574 => 209,          -- (110111.110110 | -8.15625)     => (110.10001 | -1.46875)        
    3575 => 209,          -- (110111.110111 | -8.140625)    => (110.10001 | -1.46875)        
    3576 => 209,          -- (110111.111000 | -8.125)       => (110.10001 | -1.46875)        
    3577 => 209,          -- (110111.111001 | -8.109375)    => (110.10001 | -1.46875)        
    3578 => 209,          -- (110111.111010 | -8.09375)     => (110.10001 | -1.46875)        
    3579 => 209,          -- (110111.111011 | -8.078125)    => (110.10001 | -1.46875)        
    3580 => 209,          -- (110111.111100 | -8.0625)      => (110.10001 | -1.46875)        
    3581 => 209,          -- (110111.111101 | -8.046875)    => (110.10001 | -1.46875)        
    3582 => 209,          -- (110111.111110 | -8.03125)     => (110.10001 | -1.46875)        
    3583 => 209,          -- (110111.111111 | -8.015625)    => (110.10001 | -1.46875)        
    3584 => 209,          -- (111000.000000 | -8.0)         => (110.10001 | -1.46875)        
    3585 => 209,          -- (111000.000001 | -7.984375)    => (110.10001 | -1.46875)        
    3586 => 209,          -- (111000.000010 | -7.96875)     => (110.10001 | -1.46875)        
    3587 => 209,          -- (111000.000011 | -7.953125)    => (110.10001 | -1.46875)        
    3588 => 209,          -- (111000.000100 | -7.9375)      => (110.10001 | -1.46875)        
    3589 => 209,          -- (111000.000101 | -7.921875)    => (110.10001 | -1.46875)        
    3590 => 209,          -- (111000.000110 | -7.90625)     => (110.10001 | -1.46875)        
    3591 => 209,          -- (111000.000111 | -7.890625)    => (110.10001 | -1.46875)        
    3592 => 209,          -- (111000.001000 | -7.875)       => (110.10001 | -1.46875)        
    3593 => 209,          -- (111000.001001 | -7.859375)    => (110.10001 | -1.46875)        
    3594 => 209,          -- (111000.001010 | -7.84375)     => (110.10001 | -1.46875)        
    3595 => 209,          -- (111000.001011 | -7.828125)    => (110.10001 | -1.46875)        
    3596 => 209,          -- (111000.001100 | -7.8125)      => (110.10001 | -1.46875)        
    3597 => 209,          -- (111000.001101 | -7.796875)    => (110.10001 | -1.46875)        
    3598 => 209,          -- (111000.001110 | -7.78125)     => (110.10001 | -1.46875)        
    3599 => 209,          -- (111000.001111 | -7.765625)    => (110.10001 | -1.46875)        
    3600 => 209,          -- (111000.010000 | -7.75)        => (110.10001 | -1.46875)        
    3601 => 209,          -- (111000.010001 | -7.734375)    => (110.10001 | -1.46875)        
    3602 => 209,          -- (111000.010010 | -7.71875)     => (110.10001 | -1.46875)        
    3603 => 209,          -- (111000.010011 | -7.703125)    => (110.10001 | -1.46875)        
    3604 => 209,          -- (111000.010100 | -7.6875)      => (110.10001 | -1.46875)        
    3605 => 209,          -- (111000.010101 | -7.671875)    => (110.10001 | -1.46875)        
    3606 => 209,          -- (111000.010110 | -7.65625)     => (110.10001 | -1.46875)        
    3607 => 209,          -- (111000.010111 | -7.640625)    => (110.10001 | -1.46875)        
    3608 => 209,          -- (111000.011000 | -7.625)       => (110.10001 | -1.46875)        
    3609 => 209,          -- (111000.011001 | -7.609375)    => (110.10001 | -1.46875)        
    3610 => 209,          -- (111000.011010 | -7.59375)     => (110.10001 | -1.46875)        
    3611 => 209,          -- (111000.011011 | -7.578125)    => (110.10001 | -1.46875)        
    3612 => 209,          -- (111000.011100 | -7.5625)      => (110.10001 | -1.46875)        
    3613 => 209,          -- (111000.011101 | -7.546875)    => (110.10001 | -1.46875)        
    3614 => 209,          -- (111000.011110 | -7.53125)     => (110.10001 | -1.46875)        
    3615 => 209,          -- (111000.011111 | -7.515625)    => (110.10001 | -1.46875)        
    3616 => 209,          -- (111000.100000 | -7.5)         => (110.10001 | -1.46875)        
    3617 => 209,          -- (111000.100001 | -7.484375)    => (110.10001 | -1.46875)        
    3618 => 209,          -- (111000.100010 | -7.46875)     => (110.10001 | -1.46875)        
    3619 => 210,          -- (111000.100011 | -7.453125)    => (110.10010 | -1.4375)         
    3620 => 210,          -- (111000.100100 | -7.4375)      => (110.10010 | -1.4375)         
    3621 => 210,          -- (111000.100101 | -7.421875)    => (110.10010 | -1.4375)         
    3622 => 210,          -- (111000.100110 | -7.40625)     => (110.10010 | -1.4375)         
    3623 => 210,          -- (111000.100111 | -7.390625)    => (110.10010 | -1.4375)         
    3624 => 210,          -- (111000.101000 | -7.375)       => (110.10010 | -1.4375)         
    3625 => 210,          -- (111000.101001 | -7.359375)    => (110.10010 | -1.4375)         
    3626 => 210,          -- (111000.101010 | -7.34375)     => (110.10010 | -1.4375)         
    3627 => 210,          -- (111000.101011 | -7.328125)    => (110.10010 | -1.4375)         
    3628 => 210,          -- (111000.101100 | -7.3125)      => (110.10010 | -1.4375)         
    3629 => 210,          -- (111000.101101 | -7.296875)    => (110.10010 | -1.4375)         
    3630 => 210,          -- (111000.101110 | -7.28125)     => (110.10010 | -1.4375)         
    3631 => 210,          -- (111000.101111 | -7.265625)    => (110.10010 | -1.4375)         
    3632 => 210,          -- (111000.110000 | -7.25)        => (110.10010 | -1.4375)         
    3633 => 210,          -- (111000.110001 | -7.234375)    => (110.10010 | -1.4375)         
    3634 => 210,          -- (111000.110010 | -7.21875)     => (110.10010 | -1.4375)         
    3635 => 210,          -- (111000.110011 | -7.203125)    => (110.10010 | -1.4375)         
    3636 => 210,          -- (111000.110100 | -7.1875)      => (110.10010 | -1.4375)         
    3637 => 210,          -- (111000.110101 | -7.171875)    => (110.10010 | -1.4375)         
    3638 => 210,          -- (111000.110110 | -7.15625)     => (110.10010 | -1.4375)         
    3639 => 210,          -- (111000.110111 | -7.140625)    => (110.10010 | -1.4375)         
    3640 => 210,          -- (111000.111000 | -7.125)       => (110.10010 | -1.4375)         
    3641 => 210,          -- (111000.111001 | -7.109375)    => (110.10010 | -1.4375)         
    3642 => 210,          -- (111000.111010 | -7.09375)     => (110.10010 | -1.4375)         
    3643 => 210,          -- (111000.111011 | -7.078125)    => (110.10010 | -1.4375)         
    3644 => 210,          -- (111000.111100 | -7.0625)      => (110.10010 | -1.4375)         
    3645 => 210,          -- (111000.111101 | -7.046875)    => (110.10010 | -1.4375)         
    3646 => 210,          -- (111000.111110 | -7.03125)     => (110.10010 | -1.4375)         
    3647 => 210,          -- (111000.111111 | -7.015625)    => (110.10010 | -1.4375)         
    3648 => 210,          -- (111001.000000 | -7.0)         => (110.10010 | -1.4375)         
    3649 => 210,          -- (111001.000001 | -6.984375)    => (110.10010 | -1.4375)         
    3650 => 210,          -- (111001.000010 | -6.96875)     => (110.10010 | -1.4375)         
    3651 => 210,          -- (111001.000011 | -6.953125)    => (110.10010 | -1.4375)         
    3652 => 210,          -- (111001.000100 | -6.9375)      => (110.10010 | -1.4375)         
    3653 => 210,          -- (111001.000101 | -6.921875)    => (110.10010 | -1.4375)         
    3654 => 210,          -- (111001.000110 | -6.90625)     => (110.10010 | -1.4375)         
    3655 => 210,          -- (111001.000111 | -6.890625)    => (110.10010 | -1.4375)         
    3656 => 210,          -- (111001.001000 | -6.875)       => (110.10010 | -1.4375)         
    3657 => 210,          -- (111001.001001 | -6.859375)    => (110.10010 | -1.4375)         
    3658 => 210,          -- (111001.001010 | -6.84375)     => (110.10010 | -1.4375)         
    3659 => 210,          -- (111001.001011 | -6.828125)    => (110.10010 | -1.4375)         
    3660 => 210,          -- (111001.001100 | -6.8125)      => (110.10010 | -1.4375)         
    3661 => 210,          -- (111001.001101 | -6.796875)    => (110.10010 | -1.4375)         
    3662 => 210,          -- (111001.001110 | -6.78125)     => (110.10010 | -1.4375)         
    3663 => 210,          -- (111001.001111 | -6.765625)    => (110.10010 | -1.4375)         
    3664 => 210,          -- (111001.010000 | -6.75)        => (110.10010 | -1.4375)         
    3665 => 210,          -- (111001.010001 | -6.734375)    => (110.10010 | -1.4375)         
    3666 => 210,          -- (111001.010010 | -6.71875)     => (110.10010 | -1.4375)         
    3667 => 210,          -- (111001.010011 | -6.703125)    => (110.10010 | -1.4375)         
    3668 => 210,          -- (111001.010100 | -6.6875)      => (110.10010 | -1.4375)         
    3669 => 210,          -- (111001.010101 | -6.671875)    => (110.10010 | -1.4375)         
    3670 => 210,          -- (111001.010110 | -6.65625)     => (110.10010 | -1.4375)         
    3671 => 210,          -- (111001.010111 | -6.640625)    => (110.10010 | -1.4375)         
    3672 => 210,          -- (111001.011000 | -6.625)       => (110.10010 | -1.4375)         
    3673 => 210,          -- (111001.011001 | -6.609375)    => (110.10010 | -1.4375)         
    3674 => 210,          -- (111001.011010 | -6.59375)     => (110.10010 | -1.4375)         
    3675 => 210,          -- (111001.011011 | -6.578125)    => (110.10010 | -1.4375)         
    3676 => 210,          -- (111001.011100 | -6.5625)      => (110.10010 | -1.4375)         
    3677 => 210,          -- (111001.011101 | -6.546875)    => (110.10010 | -1.4375)         
    3678 => 210,          -- (111001.011110 | -6.53125)     => (110.10010 | -1.4375)         
    3679 => 210,          -- (111001.011111 | -6.515625)    => (110.10010 | -1.4375)         
    3680 => 210,          -- (111001.100000 | -6.5)         => (110.10010 | -1.4375)         
    3681 => 210,          -- (111001.100001 | -6.484375)    => (110.10010 | -1.4375)         
    3682 => 210,          -- (111001.100010 | -6.46875)     => (110.10010 | -1.4375)         
    3683 => 210,          -- (111001.100011 | -6.453125)    => (110.10010 | -1.4375)         
    3684 => 210,          -- (111001.100100 | -6.4375)      => (110.10010 | -1.4375)         
    3685 => 210,          -- (111001.100101 | -6.421875)    => (110.10010 | -1.4375)         
    3686 => 210,          -- (111001.100110 | -6.40625)     => (110.10010 | -1.4375)         
    3687 => 210,          -- (111001.100111 | -6.390625)    => (110.10010 | -1.4375)         
    3688 => 210,          -- (111001.101000 | -6.375)       => (110.10010 | -1.4375)         
    3689 => 210,          -- (111001.101001 | -6.359375)    => (110.10010 | -1.4375)         
    3690 => 210,          -- (111001.101010 | -6.34375)     => (110.10010 | -1.4375)         
    3691 => 210,          -- (111001.101011 | -6.328125)    => (110.10010 | -1.4375)         
    3692 => 210,          -- (111001.101100 | -6.3125)      => (110.10010 | -1.4375)         
    3693 => 210,          -- (111001.101101 | -6.296875)    => (110.10010 | -1.4375)         
    3694 => 210,          -- (111001.101110 | -6.28125)     => (110.10010 | -1.4375)         
    3695 => 210,          -- (111001.101111 | -6.265625)    => (110.10010 | -1.4375)         
    3696 => 210,          -- (111001.110000 | -6.25)        => (110.10010 | -1.4375)         
    3697 => 210,          -- (111001.110001 | -6.234375)    => (110.10010 | -1.4375)         
    3698 => 210,          -- (111001.110010 | -6.21875)     => (110.10010 | -1.4375)         
    3699 => 210,          -- (111001.110011 | -6.203125)    => (110.10010 | -1.4375)         
    3700 => 210,          -- (111001.110100 | -6.1875)      => (110.10010 | -1.4375)         
    3701 => 210,          -- (111001.110101 | -6.171875)    => (110.10010 | -1.4375)         
    3702 => 210,          -- (111001.110110 | -6.15625)     => (110.10010 | -1.4375)         
    3703 => 210,          -- (111001.110111 | -6.140625)    => (110.10010 | -1.4375)         
    3704 => 210,          -- (111001.111000 | -6.125)       => (110.10010 | -1.4375)         
    3705 => 210,          -- (111001.111001 | -6.109375)    => (110.10010 | -1.4375)         
    3706 => 210,          -- (111001.111010 | -6.09375)     => (110.10010 | -1.4375)         
    3707 => 210,          -- (111001.111011 | -6.078125)    => (110.10010 | -1.4375)         
    3708 => 210,          -- (111001.111100 | -6.0625)      => (110.10010 | -1.4375)         
    3709 => 210,          -- (111001.111101 | -6.046875)    => (110.10010 | -1.4375)         
    3710 => 210,          -- (111001.111110 | -6.03125)     => (110.10010 | -1.4375)         
    3711 => 211,          -- (111001.111111 | -6.015625)    => (110.10011 | -1.40625)        
    3712 => 211,          -- (111010.000000 | -6.0)         => (110.10011 | -1.40625)        
    3713 => 211,          -- (111010.000001 | -5.984375)    => (110.10011 | -1.40625)        
    3714 => 211,          -- (111010.000010 | -5.96875)     => (110.10011 | -1.40625)        
    3715 => 211,          -- (111010.000011 | -5.953125)    => (110.10011 | -1.40625)        
    3716 => 211,          -- (111010.000100 | -5.9375)      => (110.10011 | -1.40625)        
    3717 => 211,          -- (111010.000101 | -5.921875)    => (110.10011 | -1.40625)        
    3718 => 211,          -- (111010.000110 | -5.90625)     => (110.10011 | -1.40625)        
    3719 => 211,          -- (111010.000111 | -5.890625)    => (110.10011 | -1.40625)        
    3720 => 211,          -- (111010.001000 | -5.875)       => (110.10011 | -1.40625)        
    3721 => 211,          -- (111010.001001 | -5.859375)    => (110.10011 | -1.40625)        
    3722 => 211,          -- (111010.001010 | -5.84375)     => (110.10011 | -1.40625)        
    3723 => 211,          -- (111010.001011 | -5.828125)    => (110.10011 | -1.40625)        
    3724 => 211,          -- (111010.001100 | -5.8125)      => (110.10011 | -1.40625)        
    3725 => 211,          -- (111010.001101 | -5.796875)    => (110.10011 | -1.40625)        
    3726 => 211,          -- (111010.001110 | -5.78125)     => (110.10011 | -1.40625)        
    3727 => 211,          -- (111010.001111 | -5.765625)    => (110.10011 | -1.40625)        
    3728 => 211,          -- (111010.010000 | -5.75)        => (110.10011 | -1.40625)        
    3729 => 211,          -- (111010.010001 | -5.734375)    => (110.10011 | -1.40625)        
    3730 => 211,          -- (111010.010010 | -5.71875)     => (110.10011 | -1.40625)        
    3731 => 211,          -- (111010.010011 | -5.703125)    => (110.10011 | -1.40625)        
    3732 => 211,          -- (111010.010100 | -5.6875)      => (110.10011 | -1.40625)        
    3733 => 211,          -- (111010.010101 | -5.671875)    => (110.10011 | -1.40625)        
    3734 => 211,          -- (111010.010110 | -5.65625)     => (110.10011 | -1.40625)        
    3735 => 211,          -- (111010.010111 | -5.640625)    => (110.10011 | -1.40625)        
    3736 => 211,          -- (111010.011000 | -5.625)       => (110.10011 | -1.40625)        
    3737 => 211,          -- (111010.011001 | -5.609375)    => (110.10011 | -1.40625)        
    3738 => 211,          -- (111010.011010 | -5.59375)     => (110.10011 | -1.40625)        
    3739 => 211,          -- (111010.011011 | -5.578125)    => (110.10011 | -1.40625)        
    3740 => 211,          -- (111010.011100 | -5.5625)      => (110.10011 | -1.40625)        
    3741 => 211,          -- (111010.011101 | -5.546875)    => (110.10011 | -1.40625)        
    3742 => 211,          -- (111010.011110 | -5.53125)     => (110.10011 | -1.40625)        
    3743 => 211,          -- (111010.011111 | -5.515625)    => (110.10011 | -1.40625)        
    3744 => 211,          -- (111010.100000 | -5.5)         => (110.10011 | -1.40625)        
    3745 => 211,          -- (111010.100001 | -5.484375)    => (110.10011 | -1.40625)        
    3746 => 211,          -- (111010.100010 | -5.46875)     => (110.10011 | -1.40625)        
    3747 => 211,          -- (111010.100011 | -5.453125)    => (110.10011 | -1.40625)        
    3748 => 211,          -- (111010.100100 | -5.4375)      => (110.10011 | -1.40625)        
    3749 => 211,          -- (111010.100101 | -5.421875)    => (110.10011 | -1.40625)        
    3750 => 211,          -- (111010.100110 | -5.40625)     => (110.10011 | -1.40625)        
    3751 => 211,          -- (111010.100111 | -5.390625)    => (110.10011 | -1.40625)        
    3752 => 211,          -- (111010.101000 | -5.375)       => (110.10011 | -1.40625)        
    3753 => 211,          -- (111010.101001 | -5.359375)    => (110.10011 | -1.40625)        
    3754 => 211,          -- (111010.101010 | -5.34375)     => (110.10011 | -1.40625)        
    3755 => 211,          -- (111010.101011 | -5.328125)    => (110.10011 | -1.40625)        
    3756 => 211,          -- (111010.101100 | -5.3125)      => (110.10011 | -1.40625)        
    3757 => 211,          -- (111010.101101 | -5.296875)    => (110.10011 | -1.40625)        
    3758 => 211,          -- (111010.101110 | -5.28125)     => (110.10011 | -1.40625)        
    3759 => 211,          -- (111010.101111 | -5.265625)    => (110.10011 | -1.40625)        
    3760 => 211,          -- (111010.110000 | -5.25)        => (110.10011 | -1.40625)        
    3761 => 211,          -- (111010.110001 | -5.234375)    => (110.10011 | -1.40625)        
    3762 => 211,          -- (111010.110010 | -5.21875)     => (110.10011 | -1.40625)        
    3763 => 211,          -- (111010.110011 | -5.203125)    => (110.10011 | -1.40625)        
    3764 => 211,          -- (111010.110100 | -5.1875)      => (110.10011 | -1.40625)        
    3765 => 211,          -- (111010.110101 | -5.171875)    => (110.10011 | -1.40625)        
    3766 => 211,          -- (111010.110110 | -5.15625)     => (110.10011 | -1.40625)        
    3767 => 211,          -- (111010.110111 | -5.140625)    => (110.10011 | -1.40625)        
    3768 => 211,          -- (111010.111000 | -5.125)       => (110.10011 | -1.40625)        
    3769 => 211,          -- (111010.111001 | -5.109375)    => (110.10011 | -1.40625)        
    3770 => 211,          -- (111010.111010 | -5.09375)     => (110.10011 | -1.40625)        
    3771 => 211,          -- (111010.111011 | -5.078125)    => (110.10011 | -1.40625)        
    3772 => 211,          -- (111010.111100 | -5.0625)      => (110.10011 | -1.40625)        
    3773 => 211,          -- (111010.111101 | -5.046875)    => (110.10011 | -1.40625)        
    3774 => 212,          -- (111010.111110 | -5.03125)     => (110.10100 | -1.375)          
    3775 => 212,          -- (111010.111111 | -5.015625)    => (110.10100 | -1.375)          
    3776 => 212,          -- (111011.000000 | -5.0)         => (110.10100 | -1.375)          
    3777 => 212,          -- (111011.000001 | -4.984375)    => (110.10100 | -1.375)          
    3778 => 212,          -- (111011.000010 | -4.96875)     => (110.10100 | -1.375)          
    3779 => 212,          -- (111011.000011 | -4.953125)    => (110.10100 | -1.375)          
    3780 => 212,          -- (111011.000100 | -4.9375)      => (110.10100 | -1.375)          
    3781 => 212,          -- (111011.000101 | -4.921875)    => (110.10100 | -1.375)          
    3782 => 212,          -- (111011.000110 | -4.90625)     => (110.10100 | -1.375)          
    3783 => 212,          -- (111011.000111 | -4.890625)    => (110.10100 | -1.375)          
    3784 => 212,          -- (111011.001000 | -4.875)       => (110.10100 | -1.375)          
    3785 => 212,          -- (111011.001001 | -4.859375)    => (110.10100 | -1.375)          
    3786 => 212,          -- (111011.001010 | -4.84375)     => (110.10100 | -1.375)          
    3787 => 212,          -- (111011.001011 | -4.828125)    => (110.10100 | -1.375)          
    3788 => 212,          -- (111011.001100 | -4.8125)      => (110.10100 | -1.375)          
    3789 => 212,          -- (111011.001101 | -4.796875)    => (110.10100 | -1.375)          
    3790 => 212,          -- (111011.001110 | -4.78125)     => (110.10100 | -1.375)          
    3791 => 212,          -- (111011.001111 | -4.765625)    => (110.10100 | -1.375)          
    3792 => 212,          -- (111011.010000 | -4.75)        => (110.10100 | -1.375)          
    3793 => 212,          -- (111011.010001 | -4.734375)    => (110.10100 | -1.375)          
    3794 => 212,          -- (111011.010010 | -4.71875)     => (110.10100 | -1.375)          
    3795 => 212,          -- (111011.010011 | -4.703125)    => (110.10100 | -1.375)          
    3796 => 212,          -- (111011.010100 | -4.6875)      => (110.10100 | -1.375)          
    3797 => 212,          -- (111011.010101 | -4.671875)    => (110.10100 | -1.375)          
    3798 => 212,          -- (111011.010110 | -4.65625)     => (110.10100 | -1.375)          
    3799 => 212,          -- (111011.010111 | -4.640625)    => (110.10100 | -1.375)          
    3800 => 212,          -- (111011.011000 | -4.625)       => (110.10100 | -1.375)          
    3801 => 212,          -- (111011.011001 | -4.609375)    => (110.10100 | -1.375)          
    3802 => 212,          -- (111011.011010 | -4.59375)     => (110.10100 | -1.375)          
    3803 => 212,          -- (111011.011011 | -4.578125)    => (110.10100 | -1.375)          
    3804 => 212,          -- (111011.011100 | -4.5625)      => (110.10100 | -1.375)          
    3805 => 212,          -- (111011.011101 | -4.546875)    => (110.10100 | -1.375)          
    3806 => 212,          -- (111011.011110 | -4.53125)     => (110.10100 | -1.375)          
    3807 => 212,          -- (111011.011111 | -4.515625)    => (110.10100 | -1.375)          
    3808 => 212,          -- (111011.100000 | -4.5)         => (110.10100 | -1.375)          
    3809 => 212,          -- (111011.100001 | -4.484375)    => (110.10100 | -1.375)          
    3810 => 212,          -- (111011.100010 | -4.46875)     => (110.10100 | -1.375)          
    3811 => 212,          -- (111011.100011 | -4.453125)    => (110.10100 | -1.375)          
    3812 => 212,          -- (111011.100100 | -4.4375)      => (110.10100 | -1.375)          
    3813 => 212,          -- (111011.100101 | -4.421875)    => (110.10100 | -1.375)          
    3814 => 212,          -- (111011.100110 | -4.40625)     => (110.10100 | -1.375)          
    3815 => 212,          -- (111011.100111 | -4.390625)    => (110.10100 | -1.375)          
    3816 => 212,          -- (111011.101000 | -4.375)       => (110.10100 | -1.375)          
    3817 => 212,          -- (111011.101001 | -4.359375)    => (110.10100 | -1.375)          
    3818 => 212,          -- (111011.101010 | -4.34375)     => (110.10100 | -1.375)          
    3819 => 213,          -- (111011.101011 | -4.328125)    => (110.10101 | -1.34375)        
    3820 => 213,          -- (111011.101100 | -4.3125)      => (110.10101 | -1.34375)        
    3821 => 213,          -- (111011.101101 | -4.296875)    => (110.10101 | -1.34375)        
    3822 => 213,          -- (111011.101110 | -4.28125)     => (110.10101 | -1.34375)        
    3823 => 213,          -- (111011.101111 | -4.265625)    => (110.10101 | -1.34375)        
    3824 => 213,          -- (111011.110000 | -4.25)        => (110.10101 | -1.34375)        
    3825 => 213,          -- (111011.110001 | -4.234375)    => (110.10101 | -1.34375)        
    3826 => 213,          -- (111011.110010 | -4.21875)     => (110.10101 | -1.34375)        
    3827 => 213,          -- (111011.110011 | -4.203125)    => (110.10101 | -1.34375)        
    3828 => 213,          -- (111011.110100 | -4.1875)      => (110.10101 | -1.34375)        
    3829 => 213,          -- (111011.110101 | -4.171875)    => (110.10101 | -1.34375)        
    3830 => 213,          -- (111011.110110 | -4.15625)     => (110.10101 | -1.34375)        
    3831 => 213,          -- (111011.110111 | -4.140625)    => (110.10101 | -1.34375)        
    3832 => 213,          -- (111011.111000 | -4.125)       => (110.10101 | -1.34375)        
    3833 => 213,          -- (111011.111001 | -4.109375)    => (110.10101 | -1.34375)        
    3834 => 213,          -- (111011.111010 | -4.09375)     => (110.10101 | -1.34375)        
    3835 => 213,          -- (111011.111011 | -4.078125)    => (110.10101 | -1.34375)        
    3836 => 213,          -- (111011.111100 | -4.0625)      => (110.10101 | -1.34375)        
    3837 => 213,          -- (111011.111101 | -4.046875)    => (110.10101 | -1.34375)        
    3838 => 213,          -- (111011.111110 | -4.03125)     => (110.10101 | -1.34375)        
    3839 => 213,          -- (111011.111111 | -4.015625)    => (110.10101 | -1.34375)        
    3840 => 213,          -- (111100.000000 | -4.0)         => (110.10101 | -1.34375)        
    3841 => 213,          -- (111100.000001 | -3.984375)    => (110.10101 | -1.34375)        
    3842 => 213,          -- (111100.000010 | -3.96875)     => (110.10101 | -1.34375)        
    3843 => 213,          -- (111100.000011 | -3.953125)    => (110.10101 | -1.34375)        
    3844 => 213,          -- (111100.000100 | -3.9375)      => (110.10101 | -1.34375)        
    3845 => 213,          -- (111100.000101 | -3.921875)    => (110.10101 | -1.34375)        
    3846 => 213,          -- (111100.000110 | -3.90625)     => (110.10101 | -1.34375)        
    3847 => 213,          -- (111100.000111 | -3.890625)    => (110.10101 | -1.34375)        
    3848 => 213,          -- (111100.001000 | -3.875)       => (110.10101 | -1.34375)        
    3849 => 213,          -- (111100.001001 | -3.859375)    => (110.10101 | -1.34375)        
    3850 => 213,          -- (111100.001010 | -3.84375)     => (110.10101 | -1.34375)        
    3851 => 213,          -- (111100.001011 | -3.828125)    => (110.10101 | -1.34375)        
    3852 => 213,          -- (111100.001100 | -3.8125)      => (110.10101 | -1.34375)        
    3853 => 213,          -- (111100.001101 | -3.796875)    => (110.10101 | -1.34375)        
    3854 => 214,          -- (111100.001110 | -3.78125)     => (110.10110 | -1.3125)         
    3855 => 214,          -- (111100.001111 | -3.765625)    => (110.10110 | -1.3125)         
    3856 => 214,          -- (111100.010000 | -3.75)        => (110.10110 | -1.3125)         
    3857 => 214,          -- (111100.010001 | -3.734375)    => (110.10110 | -1.3125)         
    3858 => 214,          -- (111100.010010 | -3.71875)     => (110.10110 | -1.3125)         
    3859 => 214,          -- (111100.010011 | -3.703125)    => (110.10110 | -1.3125)         
    3860 => 214,          -- (111100.010100 | -3.6875)      => (110.10110 | -1.3125)         
    3861 => 214,          -- (111100.010101 | -3.671875)    => (110.10110 | -1.3125)         
    3862 => 214,          -- (111100.010110 | -3.65625)     => (110.10110 | -1.3125)         
    3863 => 214,          -- (111100.010111 | -3.640625)    => (110.10110 | -1.3125)         
    3864 => 214,          -- (111100.011000 | -3.625)       => (110.10110 | -1.3125)         
    3865 => 214,          -- (111100.011001 | -3.609375)    => (110.10110 | -1.3125)         
    3866 => 214,          -- (111100.011010 | -3.59375)     => (110.10110 | -1.3125)         
    3867 => 214,          -- (111100.011011 | -3.578125)    => (110.10110 | -1.3125)         
    3868 => 214,          -- (111100.011100 | -3.5625)      => (110.10110 | -1.3125)         
    3869 => 214,          -- (111100.011101 | -3.546875)    => (110.10110 | -1.3125)         
    3870 => 214,          -- (111100.011110 | -3.53125)     => (110.10110 | -1.3125)         
    3871 => 214,          -- (111100.011111 | -3.515625)    => (110.10110 | -1.3125)         
    3872 => 214,          -- (111100.100000 | -3.5)         => (110.10110 | -1.3125)         
    3873 => 214,          -- (111100.100001 | -3.484375)    => (110.10110 | -1.3125)         
    3874 => 214,          -- (111100.100010 | -3.46875)     => (110.10110 | -1.3125)         
    3875 => 214,          -- (111100.100011 | -3.453125)    => (110.10110 | -1.3125)         
    3876 => 214,          -- (111100.100100 | -3.4375)      => (110.10110 | -1.3125)         
    3877 => 214,          -- (111100.100101 | -3.421875)    => (110.10110 | -1.3125)         
    3878 => 214,          -- (111100.100110 | -3.40625)     => (110.10110 | -1.3125)         
    3879 => 214,          -- (111100.100111 | -3.390625)    => (110.10110 | -1.3125)         
    3880 => 214,          -- (111100.101000 | -3.375)       => (110.10110 | -1.3125)         
    3881 => 214,          -- (111100.101001 | -3.359375)    => (110.10110 | -1.3125)         
    3882 => 215,          -- (111100.101010 | -3.34375)     => (110.10111 | -1.28125)        
    3883 => 215,          -- (111100.101011 | -3.328125)    => (110.10111 | -1.28125)        
    3884 => 215,          -- (111100.101100 | -3.3125)      => (110.10111 | -1.28125)        
    3885 => 215,          -- (111100.101101 | -3.296875)    => (110.10111 | -1.28125)        
    3886 => 215,          -- (111100.101110 | -3.28125)     => (110.10111 | -1.28125)        
    3887 => 215,          -- (111100.101111 | -3.265625)    => (110.10111 | -1.28125)        
    3888 => 215,          -- (111100.110000 | -3.25)        => (110.10111 | -1.28125)        
    3889 => 215,          -- (111100.110001 | -3.234375)    => (110.10111 | -1.28125)        
    3890 => 215,          -- (111100.110010 | -3.21875)     => (110.10111 | -1.28125)        
    3891 => 215,          -- (111100.110011 | -3.203125)    => (110.10111 | -1.28125)        
    3892 => 215,          -- (111100.110100 | -3.1875)      => (110.10111 | -1.28125)        
    3893 => 215,          -- (111100.110101 | -3.171875)    => (110.10111 | -1.28125)        
    3894 => 215,          -- (111100.110110 | -3.15625)     => (110.10111 | -1.28125)        
    3895 => 215,          -- (111100.110111 | -3.140625)    => (110.10111 | -1.28125)        
    3896 => 215,          -- (111100.111000 | -3.125)       => (110.10111 | -1.28125)        
    3897 => 215,          -- (111100.111001 | -3.109375)    => (110.10111 | -1.28125)        
    3898 => 215,          -- (111100.111010 | -3.09375)     => (110.10111 | -1.28125)        
    3899 => 215,          -- (111100.111011 | -3.078125)    => (110.10111 | -1.28125)        
    3900 => 215,          -- (111100.111100 | -3.0625)      => (110.10111 | -1.28125)        
    3901 => 215,          -- (111100.111101 | -3.046875)    => (110.10111 | -1.28125)        
    3902 => 215,          -- (111100.111110 | -3.03125)     => (110.10111 | -1.28125)        
    3903 => 215,          -- (111100.111111 | -3.015625)    => (110.10111 | -1.28125)        
    3904 => 216,          -- (111101.000000 | -3.0)         => (110.11000 | -1.25)           
    3905 => 216,          -- (111101.000001 | -2.984375)    => (110.11000 | -1.25)           
    3906 => 216,          -- (111101.000010 | -2.96875)     => (110.11000 | -1.25)           
    3907 => 216,          -- (111101.000011 | -2.953125)    => (110.11000 | -1.25)           
    3908 => 216,          -- (111101.000100 | -2.9375)      => (110.11000 | -1.25)           
    3909 => 216,          -- (111101.000101 | -2.921875)    => (110.11000 | -1.25)           
    3910 => 216,          -- (111101.000110 | -2.90625)     => (110.11000 | -1.25)           
    3911 => 216,          -- (111101.000111 | -2.890625)    => (110.11000 | -1.25)           
    3912 => 216,          -- (111101.001000 | -2.875)       => (110.11000 | -1.25)           
    3913 => 216,          -- (111101.001001 | -2.859375)    => (110.11000 | -1.25)           
    3914 => 216,          -- (111101.001010 | -2.84375)     => (110.11000 | -1.25)           
    3915 => 216,          -- (111101.001011 | -2.828125)    => (110.11000 | -1.25)           
    3916 => 216,          -- (111101.001100 | -2.8125)      => (110.11000 | -1.25)           
    3917 => 216,          -- (111101.001101 | -2.796875)    => (110.11000 | -1.25)           
    3918 => 216,          -- (111101.001110 | -2.78125)     => (110.11000 | -1.25)           
    3919 => 216,          -- (111101.001111 | -2.765625)    => (110.11000 | -1.25)           
    3920 => 216,          -- (111101.010000 | -2.75)        => (110.11000 | -1.25)           
    3921 => 216,          -- (111101.010001 | -2.734375)    => (110.11000 | -1.25)           
    3922 => 217,          -- (111101.010010 | -2.71875)     => (110.11001 | -1.21875)        
    3923 => 217,          -- (111101.010011 | -2.703125)    => (110.11001 | -1.21875)        
    3924 => 217,          -- (111101.010100 | -2.6875)      => (110.11001 | -1.21875)        
    3925 => 217,          -- (111101.010101 | -2.671875)    => (110.11001 | -1.21875)        
    3926 => 217,          -- (111101.010110 | -2.65625)     => (110.11001 | -1.21875)        
    3927 => 217,          -- (111101.010111 | -2.640625)    => (110.11001 | -1.21875)        
    3928 => 217,          -- (111101.011000 | -2.625)       => (110.11001 | -1.21875)        
    3929 => 217,          -- (111101.011001 | -2.609375)    => (110.11001 | -1.21875)        
    3930 => 217,          -- (111101.011010 | -2.59375)     => (110.11001 | -1.21875)        
    3931 => 217,          -- (111101.011011 | -2.578125)    => (110.11001 | -1.21875)        
    3932 => 217,          -- (111101.011100 | -2.5625)      => (110.11001 | -1.21875)        
    3933 => 217,          -- (111101.011101 | -2.546875)    => (110.11001 | -1.21875)        
    3934 => 217,          -- (111101.011110 | -2.53125)     => (110.11001 | -1.21875)        
    3935 => 217,          -- (111101.011111 | -2.515625)    => (110.11001 | -1.21875)        
    3936 => 217,          -- (111101.100000 | -2.5)         => (110.11001 | -1.21875)        
    3937 => 217,          -- (111101.100001 | -2.484375)    => (110.11001 | -1.21875)        
    3938 => 218,          -- (111101.100010 | -2.46875)     => (110.11010 | -1.1875)         
    3939 => 218,          -- (111101.100011 | -2.453125)    => (110.11010 | -1.1875)         
    3940 => 218,          -- (111101.100100 | -2.4375)      => (110.11010 | -1.1875)         
    3941 => 218,          -- (111101.100101 | -2.421875)    => (110.11010 | -1.1875)         
    3942 => 218,          -- (111101.100110 | -2.40625)     => (110.11010 | -1.1875)         
    3943 => 218,          -- (111101.100111 | -2.390625)    => (110.11010 | -1.1875)         
    3944 => 218,          -- (111101.101000 | -2.375)       => (110.11010 | -1.1875)         
    3945 => 218,          -- (111101.101001 | -2.359375)    => (110.11010 | -1.1875)         
    3946 => 218,          -- (111101.101010 | -2.34375)     => (110.11010 | -1.1875)         
    3947 => 218,          -- (111101.101011 | -2.328125)    => (110.11010 | -1.1875)         
    3948 => 218,          -- (111101.101100 | -2.3125)      => (110.11010 | -1.1875)         
    3949 => 218,          -- (111101.101101 | -2.296875)    => (110.11010 | -1.1875)         
    3950 => 218,          -- (111101.101110 | -2.28125)     => (110.11010 | -1.1875)         
    3951 => 219,          -- (111101.101111 | -2.265625)    => (110.11011 | -1.15625)        
    3952 => 219,          -- (111101.110000 | -2.25)        => (110.11011 | -1.15625)        
    3953 => 219,          -- (111101.110001 | -2.234375)    => (110.11011 | -1.15625)        
    3954 => 219,          -- (111101.110010 | -2.21875)     => (110.11011 | -1.15625)        
    3955 => 219,          -- (111101.110011 | -2.203125)    => (110.11011 | -1.15625)        
    3956 => 219,          -- (111101.110100 | -2.1875)      => (110.11011 | -1.15625)        
    3957 => 219,          -- (111101.110101 | -2.171875)    => (110.11011 | -1.15625)        
    3958 => 219,          -- (111101.110110 | -2.15625)     => (110.11011 | -1.15625)        
    3959 => 219,          -- (111101.110111 | -2.140625)    => (110.11011 | -1.15625)        
    3960 => 219,          -- (111101.111000 | -2.125)       => (110.11011 | -1.15625)        
    3961 => 219,          -- (111101.111001 | -2.109375)    => (110.11011 | -1.15625)        
    3962 => 219,          -- (111101.111010 | -2.09375)     => (110.11011 | -1.15625)        
    3963 => 220,          -- (111101.111011 | -2.078125)    => (110.11100 | -1.125)          
    3964 => 220,          -- (111101.111100 | -2.0625)      => (110.11100 | -1.125)          
    3965 => 220,          -- (111101.111101 | -2.046875)    => (110.11100 | -1.125)          
    3966 => 220,          -- (111101.111110 | -2.03125)     => (110.11100 | -1.125)          
    3967 => 220,          -- (111101.111111 | -2.015625)    => (110.11100 | -1.125)          
    3968 => 220,          -- (111110.000000 | -2.0)         => (110.11100 | -1.125)          
    3969 => 220,          -- (111110.000001 | -1.984375)    => (110.11100 | -1.125)          
    3970 => 220,          -- (111110.000010 | -1.96875)     => (110.11100 | -1.125)          
    3971 => 220,          -- (111110.000011 | -1.953125)    => (110.11100 | -1.125)          
    3972 => 220,          -- (111110.000100 | -1.9375)      => (110.11100 | -1.125)          
    3973 => 221,          -- (111110.000101 | -1.921875)    => (110.11101 | -1.09375)        
    3974 => 221,          -- (111110.000110 | -1.90625)     => (110.11101 | -1.09375)        
    3975 => 221,          -- (111110.000111 | -1.890625)    => (110.11101 | -1.09375)        
    3976 => 221,          -- (111110.001000 | -1.875)       => (110.11101 | -1.09375)        
    3977 => 221,          -- (111110.001001 | -1.859375)    => (110.11101 | -1.09375)        
    3978 => 221,          -- (111110.001010 | -1.84375)     => (110.11101 | -1.09375)        
    3979 => 221,          -- (111110.001011 | -1.828125)    => (110.11101 | -1.09375)        
    3980 => 221,          -- (111110.001100 | -1.8125)      => (110.11101 | -1.09375)        
    3981 => 221,          -- (111110.001101 | -1.796875)    => (110.11101 | -1.09375)        
    3982 => 222,          -- (111110.001110 | -1.78125)     => (110.11110 | -1.0625)         
    3983 => 222,          -- (111110.001111 | -1.765625)    => (110.11110 | -1.0625)         
    3984 => 222,          -- (111110.010000 | -1.75)        => (110.11110 | -1.0625)         
    3985 => 222,          -- (111110.010001 | -1.734375)    => (110.11110 | -1.0625)         
    3986 => 222,          -- (111110.010010 | -1.71875)     => (110.11110 | -1.0625)         
    3987 => 222,          -- (111110.010011 | -1.703125)    => (110.11110 | -1.0625)         
    3988 => 222,          -- (111110.010100 | -1.6875)      => (110.11110 | -1.0625)         
    3989 => 222,          -- (111110.010101 | -1.671875)    => (110.11110 | -1.0625)         
    3990 => 223,          -- (111110.010110 | -1.65625)     => (110.11111 | -1.03125)        
    3991 => 223,          -- (111110.010111 | -1.640625)    => (110.11111 | -1.03125)        
    3992 => 223,          -- (111110.011000 | -1.625)       => (110.11111 | -1.03125)        
    3993 => 223,          -- (111110.011001 | -1.609375)    => (110.11111 | -1.03125)        
    3994 => 223,          -- (111110.011010 | -1.59375)     => (110.11111 | -1.03125)        
    3995 => 223,          -- (111110.011011 | -1.578125)    => (110.11111 | -1.03125)        
    3996 => 223,          -- (111110.011100 | -1.5625)      => (110.11111 | -1.03125)        
    3997 => 224,          -- (111110.011101 | -1.546875)    => (111.00000 | -1.0)            
    3998 => 224,          -- (111110.011110 | -1.53125)     => (111.00000 | -1.0)            
    3999 => 224,          -- (111110.011111 | -1.515625)    => (111.00000 | -1.0)            
    4000 => 224,          -- (111110.100000 | -1.5)         => (111.00000 | -1.0)            
    4001 => 224,          -- (111110.100001 | -1.484375)    => (111.00000 | -1.0)            
    4002 => 224,          -- (111110.100010 | -1.46875)     => (111.00000 | -1.0)            
    4003 => 225,          -- (111110.100011 | -1.453125)    => (111.00001 | -0.96875)        
    4004 => 225,          -- (111110.100100 | -1.4375)      => (111.00001 | -0.96875)        
    4005 => 225,          -- (111110.100101 | -1.421875)    => (111.00001 | -0.96875)        
    4006 => 225,          -- (111110.100110 | -1.40625)     => (111.00001 | -0.96875)        
    4007 => 225,          -- (111110.100111 | -1.390625)    => (111.00001 | -0.96875)        
    4008 => 225,          -- (111110.101000 | -1.375)       => (111.00001 | -0.96875)        
    4009 => 226,          -- (111110.101001 | -1.359375)    => (111.00010 | -0.9375)         
    4010 => 226,          -- (111110.101010 | -1.34375)     => (111.00010 | -0.9375)         
    4011 => 226,          -- (111110.101011 | -1.328125)    => (111.00010 | -0.9375)         
    4012 => 226,          -- (111110.101100 | -1.3125)      => (111.00010 | -0.9375)         
    4013 => 226,          -- (111110.101101 | -1.296875)    => (111.00010 | -0.9375)         
    4014 => 226,          -- (111110.101110 | -1.28125)     => (111.00010 | -0.9375)         
    4015 => 227,          -- (111110.101111 | -1.265625)    => (111.00011 | -0.90625)        
    4016 => 227,          -- (111110.110000 | -1.25)        => (111.00011 | -0.90625)        
    4017 => 227,          -- (111110.110001 | -1.234375)    => (111.00011 | -0.90625)        
    4018 => 227,          -- (111110.110010 | -1.21875)     => (111.00011 | -0.90625)        
    4019 => 227,          -- (111110.110011 | -1.203125)    => (111.00011 | -0.90625)        
    4020 => 228,          -- (111110.110100 | -1.1875)      => (111.00100 | -0.875)          
    4021 => 228,          -- (111110.110101 | -1.171875)    => (111.00100 | -0.875)          
    4022 => 228,          -- (111110.110110 | -1.15625)     => (111.00100 | -0.875)          
    4023 => 228,          -- (111110.110111 | -1.140625)    => (111.00100 | -0.875)          
    4024 => 228,          -- (111110.111000 | -1.125)       => (111.00100 | -0.875)          
    4025 => 229,          -- (111110.111001 | -1.109375)    => (111.00101 | -0.84375)        
    4026 => 229,          -- (111110.111010 | -1.09375)     => (111.00101 | -0.84375)        
    4027 => 229,          -- (111110.111011 | -1.078125)    => (111.00101 | -0.84375)        
    4028 => 229,          -- (111110.111100 | -1.0625)      => (111.00101 | -0.84375)        
    4029 => 230,          -- (111110.111101 | -1.046875)    => (111.00110 | -0.8125)         
    4030 => 230,          -- (111110.111110 | -1.03125)     => (111.00110 | -0.8125)         
    4031 => 230,          -- (111110.111111 | -1.015625)    => (111.00110 | -0.8125)         
    4032 => 230,          -- (111111.000000 | -1.0)         => (111.00110 | -0.8125)         
    4033 => 231,          -- (111111.000001 | -0.984375)    => (111.00111 | -0.78125)        
    4034 => 231,          -- (111111.000010 | -0.96875)     => (111.00111 | -0.78125)        
    4035 => 231,          -- (111111.000011 | -0.953125)    => (111.00111 | -0.78125)        
    4036 => 231,          -- (111111.000100 | -0.9375)      => (111.00111 | -0.78125)        
    4037 => 232,          -- (111111.000101 | -0.921875)    => (111.01000 | -0.75)           
    4038 => 232,          -- (111111.000110 | -0.90625)     => (111.01000 | -0.75)           
    4039 => 232,          -- (111111.000111 | -0.890625)    => (111.01000 | -0.75)           
    4040 => 232,          -- (111111.001000 | -0.875)       => (111.01000 | -0.75)           
    4041 => 233,          -- (111111.001001 | -0.859375)    => (111.01001 | -0.71875)        
    4042 => 233,          -- (111111.001010 | -0.84375)     => (111.01001 | -0.71875)        
    4043 => 233,          -- (111111.001011 | -0.828125)    => (111.01001 | -0.71875)        
    4044 => 234,          -- (111111.001100 | -0.8125)      => (111.01010 | -0.6875)         
    4045 => 234,          -- (111111.001101 | -0.796875)    => (111.01010 | -0.6875)         
    4046 => 234,          -- (111111.001110 | -0.78125)     => (111.01010 | -0.6875)         
    4047 => 235,          -- (111111.001111 | -0.765625)    => (111.01011 | -0.65625)        
    4048 => 235,          -- (111111.010000 | -0.75)        => (111.01011 | -0.65625)        
    4049 => 235,          -- (111111.010001 | -0.734375)    => (111.01011 | -0.65625)        
    4050 => 236,          -- (111111.010010 | -0.71875)     => (111.01100 | -0.625)          
    4051 => 236,          -- (111111.010011 | -0.703125)    => (111.01100 | -0.625)          
    4052 => 236,          -- (111111.010100 | -0.6875)      => (111.01100 | -0.625)          
    4053 => 237,          -- (111111.010101 | -0.671875)    => (111.01101 | -0.59375)        
    4054 => 237,          -- (111111.010110 | -0.65625)     => (111.01101 | -0.59375)        
    4055 => 237,          -- (111111.010111 | -0.640625)    => (111.01101 | -0.59375)        
    4056 => 238,          -- (111111.011000 | -0.625)       => (111.01110 | -0.5625)         
    4057 => 238,          -- (111111.011001 | -0.609375)    => (111.01110 | -0.5625)         
    4058 => 238,          -- (111111.011010 | -0.59375)     => (111.01110 | -0.5625)         
    4059 => 239,          -- (111111.011011 | -0.578125)    => (111.01111 | -0.53125)        
    4060 => 239,          -- (111111.011100 | -0.5625)      => (111.01111 | -0.53125)        
    4061 => 239,          -- (111111.011101 | -0.546875)    => (111.01111 | -0.53125)        
    4062 => 240,          -- (111111.011110 | -0.53125)     => (111.10000 | -0.5)            
    4063 => 240,          -- (111111.011111 | -0.515625)    => (111.10000 | -0.5)            
    4064 => 241,          -- (111111.100000 | -0.5)         => (111.10001 | -0.46875)        
    4065 => 241,          -- (111111.100001 | -0.484375)    => (111.10001 | -0.46875)        
    4066 => 241,          -- (111111.100010 | -0.46875)     => (111.10001 | -0.46875)        
    4067 => 242,          -- (111111.100011 | -0.453125)    => (111.10010 | -0.4375)         
    4068 => 242,          -- (111111.100100 | -0.4375)      => (111.10010 | -0.4375)         
    4069 => 243,          -- (111111.100101 | -0.421875)    => (111.10011 | -0.40625)        
    4070 => 243,          -- (111111.100110 | -0.40625)     => (111.10011 | -0.40625)        
    4071 => 244,          -- (111111.100111 | -0.390625)    => (111.10100 | -0.375)          
    4072 => 244,          -- (111111.101000 | -0.375)       => (111.10100 | -0.375)          
    4073 => 244,          -- (111111.101001 | -0.359375)    => (111.10100 | -0.375)          
    4074 => 245,          -- (111111.101010 | -0.34375)     => (111.10101 | -0.34375)        
    4075 => 245,          -- (111111.101011 | -0.328125)    => (111.10101 | -0.34375)        
    4076 => 246,          -- (111111.101100 | -0.3125)      => (111.10110 | -0.3125)         
    4077 => 246,          -- (111111.101101 | -0.296875)    => (111.10110 | -0.3125)         
    4078 => 247,          -- (111111.101110 | -0.28125)     => (111.10111 | -0.28125)        
    4079 => 247,          -- (111111.101111 | -0.265625)    => (111.10111 | -0.28125)        
    4080 => 248,          -- (111111.110000 | -0.25)        => (111.11000 | -0.25)           
    4081 => 248,          -- (111111.110001 | -0.234375)    => (111.11000 | -0.25)           
    4082 => 249,          -- (111111.110010 | -0.21875)     => (111.11001 | -0.21875)        
    4083 => 249,          -- (111111.110011 | -0.203125)    => (111.11001 | -0.21875)        
    4084 => 250,          -- (111111.110100 | -0.1875)      => (111.11010 | -0.1875)         
    4085 => 250,          -- (111111.110101 | -0.171875)    => (111.11010 | -0.1875)         
    4086 => 251,          -- (111111.110110 | -0.15625)     => (111.11011 | -0.15625)        
    4087 => 251,          -- (111111.110111 | -0.140625)    => (111.11011 | -0.15625)        
    4088 => 252,          -- (111111.111000 | -0.125)       => (111.11100 | -0.125)          
    4089 => 252,          -- (111111.111001 | -0.109375)    => (111.11100 | -0.125)          
    4090 => 253,          -- (111111.111010 | -0.09375)     => (111.11101 | -0.09375)        
    4091 => 253,          -- (111111.111011 | -0.078125)    => (111.11101 | -0.09375)        
    4092 => 254,          -- (111111.111100 | -0.0625)      => (111.11110 | -0.0625)         
    4093 => 254,          -- (111111.111101 | -0.046875)    => (111.11110 | -0.0625)         
    4094 => 255,          -- (111111.111110 | -0.03125)     => (111.11111 | -0.03125)        
    4095 => 255           -- (111111.111111 | -0.015625)    => (111.11111 | -0.03125)        
  );

begin
  atan_out <= std_logic_vector(to_unsigned(LUT(to_integer(unsigned(address))),8));
end architecture;
